module lai246_290(pixels);
	//246*290
	output reg [246*290-1:0] pixels;
	always
	begin
		pixels[001*246-1:000*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[002*246-1:001*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[003*246-1:002*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[004*246-1:003*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[005*246-1:004*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[006*246-1:005*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[007*246-1:006*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[008*246-1:007*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[009*246-1:008*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[010*246-1:009*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[011*246-1:010*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[012*246-1:011*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[013*246-1:012*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[014*246-1:013*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[015*246-1:014*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[016*246-1:015*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[017*246-1:016*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[018*246-1:017*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[019*246-1:018*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[020*246-1:019*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[021*246-1:020*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[022*246-1:021*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[023*246-1:022*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[024*246-1:023*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[025*246-1:024*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[026*246-1:025*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[027*246-1:026*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[028*246-1:027*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[029*246-1:028*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[030*246-1:029*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[031*246-1:030*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[032*246-1:031*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[033*246-1:032*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[034*246-1:033*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[035*246-1:034*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[036*246-1:035*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[037*246-1:036*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[038*246-1:037*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[039*246-1:038*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[040*246-1:039*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101011011010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[041*246-1:040*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100100101011010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[042*246-1:041*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110101011101101010101010110101010010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[043*246-1:042*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011010110101010110101010101001010000100000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[044*246-1:043*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101011010111011110101010110101100000000000010010000010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[045*246-1:044*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100100100101110111110111010101001011010101010010101010010000000001000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[046*246-1:045*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000001011010101010101010101110110110101101010110100000000001000100010100001010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[047*246-1:046*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001001010111011111011111110101101101010101101001010100000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[048*246-1:047*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000100000001000100101011011110101110101011010110110111010110110101001000100000001001010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[049*246-1:048*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000010000101000000000010101101011111011111101111011011010110101011101010100000001000000000001010000100000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[050*246-1:049*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000010100100000000001001101111011110101111010111010110110101101011110011010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[051*246-1:050*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000100010000000000000011011010110101111101111101111101101111011100010100101010001000000100100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[052*246-1:051*246]=246'b000000000000000000000000000000000000000000000000000000000000000000010010100100000010010101101111111111101111110111010110111010101011101111010101000000010000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[053*246-1:052*246]=246'b000000000000000000000000000000000000000000000000000000000000000001001001000000100000000110110101010110111111011111111111010111111101011010110100100010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[054*246-1:053*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000010010000001000011101111111111111101101111101010101111010101010110101010101000000000001010000010010000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[055*246-1:054*246]=246'b000000000000000000000000000000000000000000000000000000000000000100101000000000000001101011010101011011111111101111111110101110110111001010101010101000000100000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[056*246-1:055*246]=246'b000000000000000000000000000000000000000000000000000000000000000010000100000100000000110111111111111111111111111011010111110101011010110111010101010000100000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[057*246-1:056*246]=246'b000000000000000000000000000000000000000000000000000000000000001000010000100000000101011101010101101111111111111101111010101111101101101101011010101010000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[058*246-1:057*246]=246'b000000000000000000000000000000000000000000000000000000000000100010100010000000100010111011111111111110111111111111101111011001011011011010110101010000010010100000101000001000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[059*246-1:058*246]=246'b000000000000000000000000000000000000000000000000000000000000000000001000001000000101101110101110111111111101111111011010110111101101010101001010101010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[060*246-1:059*246]=246'b000000000000000000000000000000000000000000000000000000000000001001000000000000000110110111110111111111111111110111111101111010110110101010101010000101000000001010000000100100000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[061*246-1:060*246]=246'b000000000000000000000000000000000000000000000000000000000001000000100001000000010011011101011101110111111111111101110110101101101101111011010100111000010100100000000100000001000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[062*246-1:061*246]=246'b000000000000000000000000000000000000000000000000000000000000000000001000000001000110111011111111111111111111111111101111011011011011000110010101000101000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[063*246-1:062*246]=246'b000000000000000000000000000000000000000000000000000000000000010010000000001000011101101110101011011111101111111111011010110110110100111001101001010000000001001001000001001001000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[064*246-1:063*246]=246'b000000000000000000000000000000000000000000000000000000000010000000000010000000001011110111111111111111111111011101111111101111010111010110010100101010101000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[065*246-1:064*246]=246'b000000000000000000000000000000000000000000000000000000000000001000101000100100101101011010101101111111111111111111111010110101111010101001101010010000000000000010001000000100100000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[066*246-1:065*246]=246'b000000000000000000000000000000000000000000000000000000000101000010000000000001001010110111111011111011111101110111010111101111010101101010000100100010010001001000100010000000100000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[067*246-1:066*246]=246'b000000000000000000000000000000000000000000000000000000000000000000001010000000011111101101011110111111101111111101111101011010101010010101101001010100100100000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[068*246-1:067*246]=246'b000000000000000000000000000000000000000000000000000000000000100001000000101001010101011011101011101110111110101110101111101101110111010100010100100000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[069*246-1:068*246]=246'b000000000000000000000000000000000000000000000000000000000010010100100000000000111011101110111110111111111011111011111010111011001000101010100001001010010000100010000000100100010000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[070*246-1:069*246]=246'b000000000000000000000000000000000000000000000000000000001000000000001010100001010110110101101011101011010101010110100101010110110111010001010110010000000010000000100100000000111000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[071*246-1:070*246]=246'b000000000000000000000000000000000000000000000000000000000010000000000000001010101101101111011110111101111111011101111011101101010100100100001001000001001000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[072*246-1:071*246]=246'b000000000000000000000000000000000000000000000000000000001001000100000000100001010110110101101011010110101010101010101100110101010010010010100100101000000000000100000000000000110000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[073*246-1:072*246]=246'b000000000000000000000000000000000000000000000000000000000100000000100100000010111011011110110110111101110101110111101011010101010101001001001010000100100101010000000000001000101000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[074*246-1:073*246]=246'b000000000000000000000000000000000000000000000000000000001000010000000000010100110110110101101101101011001111101100011010101010101000010010010001010000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[075*246-1:074*246]=246'b000000000000000000000000000000000000000000000000000000000010000000000010000011101101101110111011010101110010011011100101010101010010100100101010000010001001010000100000000000010000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[076*246-1:075*246]=246'b000000000000000000000000000000000000000000000000000000000100000010001000010001010110110111010101101110011101101101011010101010101001010010000101010000100000100010000000000010000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[077*246-1:076*246]=246'b000000000000000000000000000000000000000000000000000000000000100000000000001010111011011101101111011001101010101010101101010101001010001000110000000100000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[078*246-1:077*246]=246'b000000000000000000000000000000000000000000000000000000000010001000100000100101010110101011011010110111010111110101101010111011010101010011000101010001000000010000001000000000100000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[079*246-1:078*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000100000011101101111101110101101110111101011110110111001101010100101000101000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[080*246-1:079*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000001001010110110101010111110111011110110101011011010110110110110010110100101001010000101000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[081*246-1:080*246]=246'b000000000000000000000000000000000000000000000000000000000001010010010000000010101011011111101011101111011011111101010111111011101010101001010000100000000000000001000001000010000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[082*246-1:081*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000100001011011110110101011110111011111110101011101110101110010101001010001010001000101000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[083*246-1:082*246]=246'b000000000000000000000000000000000000000000000000000000000001000000000000100101101001101111111011111110110111110110111011111101110101010101010000100010000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[084*246-1:083*246]=246'b000000000000000000000000000000000000000000000000000000000000001001000000001010110110110101011111010111111101011011011101110110101010101000101010001000000010000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[085*246-1:084*246]=246'b000000000000000000000000000000000000000000000000000000000000100000000100100111011011011111110101111011010111101110110111011011010101010101000001000001010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[086*246-1:085*246]=246'b000000000000000000000000000000000000000000000000000000000000000000010000001010110110101010101111101110111101010101101010110110101010101010101010000100000000001000000000010101000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[087*246-1:086*246]=246'b000000000000000000000000000000000000000000000000000000000001001000000000101101101101111101111010111011101011111011011101101001010101010101010100101000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[088*246-1:087*246]=246'b000000000000000000000000000000000000000000000000000000000000000001000010000110110111010111011111101101010101010101101010110110101010101010101010000010100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[089*246-1:088*246]=246'b000000000000000000000000000000000000000000000000000000000000100000000000101011011101101101101010110110111010101111010110101001001010101010010010101000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[090*246-1:089*246]=246'b000000000000000000000000000000000000000000000000000000000000001000000000001110111011011011011111101101100101011000110101010101010101010100100100100001001010010000000100010000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[091*246-1:090*246]=246'b000000000000000000000000000000000000000000000000000000000001000000010001010101101110110110110101011011011010100111001010101010101000101010101010010100010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[092*246-1:091*246]=246'b000000000000000000000000000000000000000000000000000000000000000010000000011010110101011011011010101101001010110101101001010101010110010001010001000010000010000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[093*246-1:092*246]=246'b000000000000000000000000000000000000000000000000000000000000101000000001001111011011101101101111010010110001001010010010000000000001000110000100101001001000100000000000010100000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[094*246-1:093*246]=246'b000000000000000000000000000000000000000000000000000000000000000000001000011010110111011011010101010101001010010100100100010101010010011000101001000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[095*246-1:094*246]=246'b000000000000000000000000000000000000000000000000000000000000000010000000101111101100110110111010100000010000101010001001000000000101000110100010010100101000000100001001010000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[096*246-1:095*246]=246'b000000000000000000000000000000000000000000000000000000000000010000100000010101010111011011010101010101001010010101000100101011101000110001011000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[097*246-1:096*246]=246'b000000000000000000000000000000000000000000000000000000000000001000000010011011111010101101111010001000010001000000010010000010000010001010100101010101001000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[098*246-1:097*246]=246'b000000000000000000000000000000000000000000000000000000000000000001010000100111010110111011010101010010100010011111100000110100010101010100001010000000010010100000100010100000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[099*246-1:098*246]=246'b000000000000000000000000000000000000000000000000000000000000001000000000101111110101001010101010100100010100101100010101001001000000001001010000101010000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[100*246-1:099*246]=246'b000000000000000000000000000000000000000000000000000000000000000010100100110101011010110101010101010010001010000010001000100100101010100100001010010001010101000100001000100000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[101*246-1:100*246]=246'b000000000000000000000000000000000000000000000000000000000000000000010001010111010110101010000000000100100001010100100010010010000000000000100001001100101000100000100010000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[102*246-1:101*246]=246'b000000000000000000000000000000000000000000000000000000000000000101000100011010101100100000101010101001010111000101000100100000100100000010000010010101000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[103*246-1:102*246]=246'b000000000000000000000000000000000000000000000000000000000000000000010001101011010111010100000000000010000100011011010010101010000001010100100100111000010000100001001010000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[104*246-1:103*246]=246'b000000000000000000000000000000000000000000000000000000000000000001000100110101110101001011010101010001010011001110101001000000101000000010010000001101000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[105*246-1:104*246]=246'b000000000000000000000000000000000000000000000000000000000000000000100001011110101111111101101000100100001000010111110100101010000010101001001010100000010001010000100100000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[106*246-1:105*246]=246'b000000000000000000000000000000000000000000000000000000000000000001000100110101111010100101011011001001010011010101101001000000010100000010010000000101000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[107*246-1:106*246]=246'b000000000000000000000000000000000000000000000000000000000000000000010001011010110111111010100100010010000100101111011101010101000001010100100101010000001001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[108*246-1:107*246]=246'b000000000000000000000000000000000000000000000000000000000000000000100100101111011110110101010010101001110101001111100100000000101000000010010000001001000000100000101000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[109*246-1:108*246]=246'b000000000000000000000000000000000000000000000000000000000000000000010001011010111111111110100100000010011010010110111010110101010010101001000101010100001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[110*246-1:109*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000100110111101011011111101001111111111111011111110101001010000101010010001010100000010000101000010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[111*246-1:110*246]=246'b000000000000000000000000000000000000000000000000000000000000000000010001011101011111111011111111011111111010111111011010101111110010001001010011001010100101000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[112*246-1:111*246]=246'b000000000000000000000000000000000000000000000000000000000000000000001000101111100101111111111111111111101001010111101101100001011001101101011100100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[113*246-1:112*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000100101010110111011111011011111101110100111110111010010101101110110110101010010010010101010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[114*246-1:113*246]=246'b000000000000000000000000000000000000000000000000000000000000000000001001011101101011111111111111101011010101101111010010100010111101101101110100100100100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[115*246-1:114*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000010100111010110111111110101010100001011111111101100001001010111111011010101001000001010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[116*246-1:115*246]=246'b000000000000000000000000000000000000000000000000000000000000000000001000011011111011010101011010101010100010101101110010100000001001011101101101100101000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[117*246-1:116*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000101010110101101101010100101010001001011110111010100011101010010101010111010010000010100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[118*246-1:117*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000010011010111011110100101010100010011111011101010001101000000101001010100111010010100000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[119*246-1:118*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000100101101101110101001001001001000110101110110100110110110010000010101011000100100001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[120*246-1:119*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000011010110110111110100100100100101011110101011010001011001000101001010101110010001000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[121*246-1:120*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000101010101011010101010010010010000111111011100101010100100010000100100000001000100010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[122*246-1:121*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000011010101110101101000100100000101110010101011000000001000000101001000101010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[123*246-1:122*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000010101010101110010101001001010001001101010100010101010010100000010010010100100010001010010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[124*246-1:123*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000111010110110011101000100100000100100101010010100000001000001001001001000010010001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[125*246-1:124*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000010101101001100101010010000100010010000100100001010100010000100000100101001000100010100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[126*246-1:125*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000110101010110101010000100010000100100010001001010000000000010000010001000010001010100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[127*246-1:126*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000101010101010100101001000101001000100000010000010001000100010100100010100100000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[128*246-1:127*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000010101010101010010100100000100010001010000001000100010001000000010000010010101010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[129*246-1:128*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000001010101010001000010010010001010000000000100000000000000000101000101000100010000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[130*246-1:129*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000010101010101010010100000000100110010000010000010001000100010000001010001000100101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[131*246-1:130*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000001010101000101000001001001011011000101000001000000010001000010100000100101001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[132*246-1:131*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000001101010110000101000100000001101111010000100001000000000001000010101010010100101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[133*246-1:132*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000010101001101010010010010110110101010100000100001001010000001000000001000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[134*246-1:133*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000101010010010000100000000101101010001000010000100000000100100010101010010100010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[135*246-1:134*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000010101101001010001010101010010000100010000010000101001000000100000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[136*246-1:135*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000011010100100101000000000001001010010001010000100000100010010001010100010100101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[137*246-1:136*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000101011010000010101010100100001000100001010000100001001000100001001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[138*246-1:137*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000011010100101010100000000000001010001001010000010000000000010001010010010100101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[139*246-1:138*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000101011010000001001000001000000010000000100000000000000000100000100100001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[140*246-1:139*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000010110100101101000100010000000000000000000000000001001010010001010010010100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[141*246-1:140*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000001001011010010010010000100010001000010010000100100000000000100001001000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[142*246-1:141*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000011010010100100000010001000100001000000010000000010000010001010000010100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[143*246-1:142*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000100101101010001010000100101010100001000000001000100101000100000101000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[144*246-1:143*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000110100101001100001010010100101010100010100100010000000010010100000101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[145*246-1:144*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000001011010010010100000001011000010010000000001000010010000000001010000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[146*246-1:145*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000011010010100100000010101000101000100100010100001000000100101010100101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[147*246-1:146*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000010101101010001010100010101001010001001000001000010100001000000001000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[148*246-1:147*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000010110010101000000010101010100001000000001000010000010000010101010101010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[149*246-1:148*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000001001101010101010100101010010100000100100001001010000101000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[150*246-1:149*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000010111010101000000011011010100000010000000100000000010000000100101010100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[151*246-1:150*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000010100101010010101101100101010010100101001001010010000100101001000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[152*246-1:151*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000001011010101001010100111110101000000000000000001000100010000100100010100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[153*246-1:152*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000101010111010110001011010011010101010100100101000010010000010010001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[154*246-1:153*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000000010110100101001010110101110110110000000000000001000000010100100010010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[155*246-1:154*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000001101010111010110101001110101011001010010101001000010101000001001000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[156*246-1:155*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000010111101010111010010110011010101010001000000000010000000101000000100010010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[157*246-1:156*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000000101011110101100101010101100101010100100100100101000101010000101010001001000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[158*246-1:157*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000001011110101101011101010101001010100001000001001000010000000010000000010000001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[159*246-1:158*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000011111111110010101010101010110100010100010100000001000101001000101010100101010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[160*246-1:159*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000000111111101011101010101010101000010001010000010101000010000100010000000010000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[161*246-1:160*246]=246'b000000000000000000000000000000000000000000000000000000000000000000000111111111111110101010110101010110100100000101000000101001010001000100101000010010001000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[162*246-1:161*246]=246'b000000000000000000000000000000000000000000000000000000000000000000011111111111101101110010101010101001001010101000010101000010000100010001000010100100100010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[163*246-1:162*246]=246'b000000000000000000000000000000000000000000000000000000000000000111111111111111011011010101010101010101010100010010100000010100100001000100010000000000001000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[164*246-1:163*246]=246'b000000000000000000000000000000000000000000000000000000000000111111111111111111111111011010101010100100101011001001010101000010010100010001001001010010000001001000101000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[165*246-1:164*246]=246'b000000000000000000000000000000000000000000000000000000000111111111111111111111101101110100010101010101010000100100001000101000000001000100000100001000100100000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[166*246-1:165*246]=246'b000000000000000000000000000000000000000000000000000000111111111111111111111111111110101101101010101010100101001001010101000010100100010001010000100010000000010000110101010000000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[167*246-1:166*246]=246'b000000000000000000000000000000000000000000000000000111111111111111111111111111111011101010000010101010010010010010100000010100001001000100000101001000010010000100001010101010000000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[168*246-1:167*246]=246'b000000000000000000000000000000000000000000000000111111111111111111111111111111111110111010110100010101011001001000010101000010100000010001010000000010000000100001010001001001010000000000000000000000000000000000000000000000000000000000000000000000;
		pixels[169*246-1:168*246]=246'b000000000000000000000000000000000000000000000111111111111111111111111111111111111111101101001010100010100110110011001010101000000101000100000010101000100100010000001010100110101010000000000000000000000000000000000000000000000000000000000000000000;
		pixels[170*246-1:169*246]=246'b000000000000000000000000000000000000000001111111111111111111111111111111111111111011011010010001010101001001000100010000000010010000010000100100000000000001000101010101001001010101010000000000000000000000000000000000000000000000000000000000000000;
		pixels[171*246-1:170*246]=246'b000000000000000000000000000000000000101111111111111111111111111111111111111111111110110111010100001000100100101010100101010100100100100100001000100101001000000000010010100100101010101010000000000000000000000000000000000000000000000000000000000000;
		pixels[172*246-1:171*246]=246'b000000000000000000000000000000000111111111111111111111111111111111111111111111111111111010101010100100010010010000010000000000000010000010100010010000000010010001001001010110010101010101010000000000000000000000000000000000000000000000000000000000;
		pixels[173*246-1:172*246]=246'b000000000000000000000000000000111111111111111111111111111111111111111111111111111111101111010001001001001001000101001010101010101000101000001000000100010001000100101010101001100010001010101010000000000000000000000000000000000000000000000000000000;
		pixels[174*246-1:173*246]=246'b000000000000000000000000000011111111111111111111111111111111111111111111111111111101011010100110010010010010001000010000000000000010000000100001010001000100000001010010010010001100110101010110110000000000000000000000000000000000000000000000000000;
		pixels[175*246-1:174*246]=246'b000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111011001000100100100100010100101010101001000100101001000000000000000101000101001001010110010101010101001001101000000000000000000000000000000000000000000000000;
		pixels[176*246-1:175*246]=246'b000000000000000000000001111111111111111111111111111111111111111111111111111111111111101011100100110010010010010000010000000000100010010000000100100100101000000010100101101001001010010001010101100101010000000000000000000000000000000000000000000000;
		pixels[177*246-1:176*246]=246'b000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110110101001001001001000101001010101010001000001001010010010000000001001001011010000110110100100110101010011010100100000000000000000000000000000000000000000000;
		pixels[178*246-1:177*246]=246'b000000000000000000011111111111111111111111111111111111111111111111111111111111111111110101101010010010010010101000010000000000100010100010000000000010100010000010100100111001000101101001010101010010101101000000000000000000000000000000000000000000;
		pixels[179*246-1:178*246]=246'b000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111010100100100100100000101000101010100001000001000100100100000001000010101010011000101011010010110001010101101010010100000000000000000000000000000000000000000;
		pixels[180*246-1:179*246]=246'b000000000001111111111111111111111111111111111111111111111111111111111111111111111111111101111010010010010010100000100000000010100010100010010000001000100001001010001000110100100101001001100101010010101010111000000000000000000000000000000000000000;
		pixels[181*246-1:180*246]=246'b000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111101010101001001000001010001010101000001000001000001001000010000100100100110111000011011010101010011010010101010101000110000000000000000000000000000000000000;
		pixels[182*246-1:181*246]=246'b000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000010010001010000010000000000100000100000100000010000010001001001001000011100100101010010100100101010101011011101100000000000000000000000000000000000;
		pixels[183*246-1:182*246]=246'b000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010100100100000101000101010101001010001010000100000100000010110110101011010010101010101101011010101010111101101011111100000000000000000000000000000000;
		pixels[184*246-1:183*246]=246'b000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100010010010100000100000000000000000100000010001000001001001001001010100101010010101010010100101010101010110111101111111100000000000000000000000000000;
		pixels[185*246-1:184*246]=246'b000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001001001000001010010101001001010010010001000000010000100110101010101001010101101010100101011010101010111111110111111111111100000000000000000000000000;
		pixels[186*246-1:185*246]=246'b010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010010001010000000000010000000000000100010010000101001101010101010010100010010100101010100101010101101011011111011111111111000000000000000000000000;
		pixels[187*246-1:186*246]=246'b101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100100100000101010010000010010100100000000000101010110010101010001101011001101011010101011010101011011111111111111111111111110000000000000000000000;
		pixels[188*246-1:187*246]=246'b110111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111110110100010010000000000100000000000000010001010101010011001000101100010100100010100101000100101010111101111111111111111111111111110000000000000000000;
		pixels[189*246-1:188*246]=246'b011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111101100100100100000100100010101000110101010101100101011010101101011011101010101011011010101110111111111111111111111111111111100000000000000000;
		pixels[190*246-1:189*246]=246'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111010101011011001010101001001101010111010101010101001010100100010010100100010101010100010010101011111111111111111111111111111111111000000000000000;
		pixels[191*246-1:190*246]=246'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101111011010101110101110110110010101001010110101010110100101011001001010101101010101011001101101111111111111111111111111111111111111110000000000000;
		pixels[192*246-1:191*246]=246'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110101101111110101110011011011101010110101010110101010010010100101100101010010101010100110101011111111111111111111111111111111111111111100000000000;
		pixels[193*246-1:192*246]=246'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010010110101101010101011101101011010101010101101101011010011010010101010101011001010111011111111111111111111111111111111111111110000000000;
		pixels[194*246-1:193*246]=246'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011110101101101011010111011010011010110101010101010010010100010100010101010010101010010101111111111111111111111111111111111111111111110000000000;
		pixels[195*246-1:194*246]=246'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101111011011101101010101101100101001010101010001010101011001011101010101101010101101010111111111111111111111111111111111111111111100000000000;
		pixels[196*246-1:195*246]=246'b111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111010101101010101011101100110111010110101010101101001010100101000010101010010101010101011111011111111111111110111111111111111111111110000000000;
		pixels[197*246-1:196*246]=246'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111010010110101010010011001000101001010101010010110101011010111101010010101010101010101011111111111111111111111111111111111111111111000000000;
		pixels[198*246-1:197*246]=246'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101110101010101101101011011010110101010100101001010100010100010010101010101010101010111111111111111111111111111111111111111111111100000000;
		pixels[199*246-1:198*246]=246'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110101010101010101010100100101001010100101010110101011101011010101010101010101010101111111111111111111111111111111111111111111111000000000;
		pixels[200*246-1:199*246]=246'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111011011010101010101010110101101010010010101001010100010100101010101010101011011010111111111111111111111111111111111111111101111110000000;
		pixels[201*246-1:200*246]=246'b111111110111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111010110110101010101010101001010010101101101010110100101101011010101010101010110100111111110111111111111111111111111111111111111011111000000;
		pixels[202*246-1:201*246]=246'b111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101101011010101010101011010101010010010101000101001010100101010101010010101011101011111111101111111101111111111111111111010110111000000;
		pixels[203*246-1:202*246]=246'b111111011111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111101011011101101010101010100101010101010101010111010110101011010101010101101010110011111111111111111111111111111111111111111111111101100000;
		pixels[204*246-1:203*246]=246'b111101111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101010110101010101010101001010101010101000101010101001010101001010010101011101111111111111111111111111111011111111110101101111110000;
		pixels[205*246-1:204*246]=246'b111111111111110111110111111111111110111111111111111111111111111111111111111111111111111111111111111111111111110110110110101010101010101010110101010101010111010101010110101010110101101010101010111101111111111111011111111111111111111111111011110000;
		pixels[206*246-1:205*246]=246'b111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101101010111010101010101001010010101010100101001010101010101001010010101110111111111111111111111111111111111111111110111111110110000;
		pixels[207*246-1:206*246]=246'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011101001101110101010110101101010101011010110101010101010110101101010011101111111111111111111111111111111111111011110111111111000;
		pixels[208*246-1:207*246]=246'b111111111111111111111111111111110111111111101111111111111111111111111111111111111111111111111111111111111111111111101100111110110011010101010100101010101001010010101010101010010100101011101110111111110111111110111111110111111111101111101101111100;
		pixels[209*246-1:208*246]=246'b111111111111111111111111111011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111011101001001110111010101011010101010110101101010101010101101011010100010111111111111111111111101111111111111110110111111111101100;
		pixels[210*246-1:209*246]=246'b111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010110111001100101101010110101010100101001010101010101001010101011101111111111111111111111111111111111111111101101011111111100;
		pixels[211*246-1:210*246]=246'b111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011010110011110010101001010101011010110101010101010110101010100111111111111011111111110111111110111110110111111111110110110;
		pixels[212*246-1:211*246]=246'b111111010110111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111110110101101011100011101101110110110101010010101010101010010101010111001111111111111111111111011111111111111111101110111011111110;
		pixels[213*246-1:212*246]=246'b111111111011111111111101111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111101101010101011101011010101101001010101101010101010101010101010100111011111111111111111111111111111111111101111111011111011010;
		pixels[214*246-1:213*246]=246'b111101101111111111111111011111111011111111111111111111111111111111111111111111111101111011111111111111111111111111111111111011011010101011010110101010110101101010101010101010101010101011010111111111111101111111011111101111111111111011111111111110;
		pixels[215*246-1:214*246]=246'b111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111101101100101110100101011010101101010010101010101010101010101010101111111111111111111111101111111111111111011101111111110110110;
		pixels[216*246-1:215*246]=246'b111111111111110111011111111111111111111111111111111111011010110111111111101111111111111111110111111111011111111011111111110100111010010111010101010110101101101010101010101010101010101110101111101111111111111110111111111111111111111101110111111110;
		pixels[217*246-1:216*246]=246'b101101111111111111111111101111111111111111111111111101111111111111011111111111111111111111111111110111111111111111110111111111010101010100101010101001010010010101010101010001010101011001111111111111111111111111011111101111110111110111111111011010;
		pixels[218*246-1:217*246]=246'b111111011111111111111111111111111111111111111111110111101011111111110111111111101111011111111111111111110111111110111101111010101010110101010101011010110101101011010101010110100101010110111111111111101111111101111111111111111111101111111010111110;
		pixels[219*246-1:218*246]=246'b111111111111111111111110111111111111111111111101111111011111111111111111111111111111111111111111111111111111111111111111111111010101001011010101010111010101010100101010101001010101010101111111111111111111111111011111111111101111110111011111101101;
		pixels[220*246-1:219*246]=246'b111011111111111111101111111111111111111111110111011011111111111111111111111111111111111111111111111111111111111111111111111101111010110101010101101001010101010111010101001010101010101010111111111111111111011101111111011111111111011011110101110111;
		pixels[221*246-1:220*246]=246'b011111111111111101111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111010110101010101010010110101010101100101010110101010101010101111111111111111111111110111111111111111111101111111111011101;
		pixels[222*246-1:221*246]=246'b111111011011011111111111111111111111111111011101101011111111111111111111101111111111111111111111111111111111111111111111111111111101010101010101110100101101101011010110100101010100101011111111111011111011111111111111111111011111110111101010111111;
		pixels[223*246-1:222*246]=246'b111111111111111111111110111111011111111101111111011111111111111111111111111110111111111111101111111111111111011111111111111111111010101010101010001011010110010100101001011010101011010101111111111111111111111110111111111111111101011111011011101010;
		pixels[224*246-1:223*246]=246'b111010111111111111101111111111111111110111110101111111111111110111111111111111111111111011111111101111111111111110111111111111111111010101010101101100101011101011010110101010100100101011111111011111111111111111011111011110111111101111101101111101;
		pixels[225*246-1:224*246]=246'b101111011111111111111111111111111111111111011111011111111111111111111011111111111111111111111111111111011111110111111101101111111111111010101010010011010100010100101011010101011011010111111111111110111011111111111111111111110101110110111010101011;
		pixels[226*246-1:225*246]=246'b111011111111111110111111111111111111111101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111010101101010101011100101101111110101010100101010110111101011111111011110111111111111111011101111100111110110;
		pixels[227*246-1:226*246]=246'b101110111111110111101111111111111110101111010111111111111111111111011111111111101111111111111101111111111111111111111111111111111111111101011010010101001010011010010011111110101011010101101111011111111101111111111111111111101111011110111010101011;
		pixels[228*246-1:227*246]=246'b111111111111111111111111110111111111111011111111111111111111111111111111101111111111111111110111111101111111111111110111111011111111011111101101010101101011001001011101111011110100101010010101101011111111111111011111011011110111101111001111111101;
		pixels[229*246-1:228*246]=246'b110111111111110101111101111111111011101110101111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111101010010100110110100101111111111111010101101010110101111111110111111111111111010111111010101001001010;
		pixels[230*246-1:229*246]=246'b111111111111011111101111111111111110110101111111111111111111111111111111111111111111110111111111111111111111111011111111111111111111111111111110101010110101100100101011111111111110111010011101101111101110111111111111111110101111101111110110111011;
		pixels[231*246-1:230*246]=246'b111111111111110111111111111111101111011111011111111111101111101111111111111111111101111111111111111111111111111111111111111111101111111111111111111101001010011011010101111111111111111110100110101011111111111101101111111111011110111010011011010101;
		pixels[232*246-1:231*246]=246'b111111111101111011111111111111111010101011111111111111111111111111111111111111111111111111111111111111111110111111111101111111111111111111111111111110101011001001011011110111110111111111111010110101111101111111111111110101101111101101101011101101;
		pixels[233*246-1:232*246]=246'b111111111110101111011011111111101101111111111111111111111111111111011101111111111111111110111110111011111111111111011111101101111110111110111011111111110100101010100111111111111111111011011011001011011111111110111111111111011111111011010101011010;
		pixels[234*246-1:233*246]=246'b111111111111111011111111111110111011101111111111111101111101111111111111101111111111111111101111111110111111101111111111111111111111111111111111111111101101010101011111111101111111111111111110111110111011011111110111011100101111010110110110110111;
		pixels[235*246-1:234*246]=246'b111111111101101110110111111111101101111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111101111111011111111011111111010101010101111111111111111111111111111101001101110111111111111110111011111101010101011010100;
		pixels[236*246-1:235*246]=246'b111111111111010111111111111101010111111111111111111111111111111011111111111111111111111111111111111111111111111111011011101111111111111111111111111111111110101010111111101111111101111111011011111111011111111011011111111001111110110101010101101011;
		pixels[237*246-1:236*246]=246'b111101110101111010101011011111111011111111111111111111111111111111111111111111111110111111111111101111111111111111111111111111111111111111011111111101111111010101111111111111111111111111111111101101101011011111101111101111001111101110101110110110;
		pixels[238*246-1:237*246]=246'b111111111111101111111111111010101111111111111111111111111111111111111111111111111111111011111111111110111111110111111111111110110111111111111011111111111111111111111111111101111111111111111111111111011111111110111110110100111101011001011001101101;
		pixels[239*246-1:238*246]=246'b101111101010111010110111111101110111111111111111111111111111111111111111111111111111111111111011111111111111111111111101111111111111011110111111011111101111111111101111111111111110111111111101111011110101111011101111101101111111010111100110101010;
		pixels[240*246-1:239*246]=246'b111111111111011111111011110110101111111101111101111111011111111111111111111111111111111111111111111111111011111111011111101111111111111011111101110101111111101111111111111111110111111101011111011110101111011111110111110110111101101010111011010101;
		pixels[241*246-1:240*246]=246'b110110110101101010011111111011111111111111101111110111111111011111111111011111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111101111101010111010101011110110101001010111011;
		pixels[242*246-1:241*246]=246'b011111101111111101110111010101011111111111111111111111111111111101111111110111011111111111111111111111111111111111111111111111111111111111111111111111011101111111111111111111111111101111111111111101101111011011101110111010111111101110110101100110;
		pixels[243*246-1:242*246]=246'b110101111010101011011111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111101111111111111111111111111111111101101111111111111111111111111111101111111010110110110111010111011100101001011010101010;
		pixels[244*246-1:243*246]=246'b111110101111110101111101001011111111111111111111111111110111111111111111111111111110111111111111111111111111111111111111111101111111111111111111111111111111011111111111111110111111111111110101111111011101011011011101101001111111010110101101011101;
		pixels[245*246-1:244*246]=246'b101011110101011110110111110111111111111111111111111111111111111111111111111111111111111111101101111111111011110111011111111111111111111111111111111111111111111111111011111111111111011111111111111101110110101110100111011101011010101101101011101010;
		pixels[246*246-1:245*246]=246'b011111011111110101011101011111111111111101111111011101111111111111111111111111101111111111111111011111111111111111111110111111111111111011011110111111011111110111101111111111110111110111111111011011010101111001111110110010111110111011010110011011;
		pixels[247*246-1:246*246]=246'b110101110101011011110111101011111111101111111011111111111110111011111111101111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111110111011111111101010010110001010101101110101001010110101100100;
		pixels[248*246-1:247*246]=246'b111110111111101101011100111111111101111111111111111111111111111111110111111111111111011011111111111101111111111111111111111011111111111111111111111111111101111111111111111110111111111111111110101010111011101011111101110101111011110101011010111011;
		pixels[249*246-1:248*246]=246'b101011101010110101110111010111110111111111111111111111111111111111111111111111111111111111111111111111111011111111101111111111111110111111111111011111111111111111111111111011111011101111111111111111101100011101010011001011110110101011010101010110;
		pixels[250*246-1:249*246]=246'b011111011101101011101110101111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111101011111111111111111111111111111011111111011110111011110111111111111011111111010101011110010101110110010101100101110110110110101;
		pixels[251*246-1:250*246]=246'b110101110111011101011011111111101111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111110111111111110111111111111111111101111111111111111111011101111110101011101011100011101010101010111010101110101011011001010;
		pixels[252*246-1:251*246]=246'b101110101010100111101010011110111111111111011111111110111011111111111111111111111111111111110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110101111101011000110111011011010110110011011001010110101;
		pixels[253*246-1:252*246]=246'b111011111111111101010101111011111111111111111111111111111111111111111101110111111111111111111111111111111111111111111111111111111111111111111011111101111111111111111111111111011111111111011111110101010110111010101010101101101101110110110110101011;
		pixels[254*246-1:253*246]=246'b010110101010101010101011101110111111101111111111101111111111111111111111111111111110111011111111111111111111111110111111111111111111111111111111011111111011111111111111111111111111111011111010111111101001100101010101011010101011001101101101010110;
		pixels[255*246-1:254*246]=246'b111101110111010111010110110101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111110111111111111111111111111011101101111011110111111111111101111101010110110011010101010110111010101110010010010111010;
		pixels[256*246-1:255*246]=246'b101110111001101010101011011111111111111101111011111111111111111111011111111111101111111111111111111111111111011111111011111111110111111111111111111111111111111111111101111111111101101110111110111101011011010101010101011001101110011101101101001101;
		pixels[257*246-1:256*246]=246'b011011010111011101010100101010111111111111111111111111111111111111111111111111111111110111111011110111101111111111111111111111111111111111111111111111111111111111111111101111111111111011110111010111100101010101001011110110110101110011011010110011;
		pixels[258*246-1:257*246]=246'b110110111010101011101001101011111111111111111111111111111111111111111111111110111111111110101111011101111111111111111111111111111111111111111111111111111111111011111111111111111111111111111110111010011010110100010101001101101011001110101011101110;
		pixels[259*246-1:258*246]=246'b101101101101011111010110010111111111111111111111111111111111111111111111111111111110111111111010111111111101111010111011011011011111110111011111101101101111111111101111111110111011111011010111101101101101001001011010110110110101110101010101010101;
		pixels[260*246-1:259*246]=246'b110110110110101010101001011010101111111111111111111111111110111111111111011111111111111111101111101111011111011111101111111111111010111111111010111111111011111111111111011011101111011101111010110110110101110100101101011011011110011010111010110110;
		pixels[261*246-1:260*246]=246'b011011101001011110101010100101111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111001101001101101011001010010011101010101001110101100110101101;
		pixels[262*246-1:261*246]=246'b111101011110110001010101011011011111011111111111111111111111111011111111111111111111110111111111111111111111111111111101110111111111111111111111111111111111111111111111111111111101111101111010111011001010111010101101010110110111001011011101011001;
		pixels[263*246-1:262*246]=246'b101011010011001110101010101101111101111111111111110111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111011111011111010101111101010101010110101011011010110101010010101110;
		pixels[264*246-1:263*246]=246'b110110101101100010110101010110101111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111011111011011011111111111111111111101101101111111011111110111101010101100100110101010111011011101101011011110101101110011;
		pixels[265*246-1:264*246]=246'b011101101011011101001010101010111111111111111111111111111111111111111111111011111101111111111111111011111111111101111111111111111111111111111111111110111111111111111111111011110110111010111101111011010101101001001010110010101100101001011010101010;
		pixels[266*246-1:265*246]=246'b101011010110101010110101010101011111111111011101111111111111111111111111111111011111011110110110111111111111011111011111111111111011111111111101110111111101111111111111101111111111101111101011000110111101010010110110101111011011110110110111101101;
		pixels[267*246-1:266*246]=246'b111010111001010101010100101111111111111011111111111111111111111111111111111111111111111111111111111111011111111111111111011111111111111111111111111111111111111111111011011101011011111010110101111011010110101001011010101001100101001011010100110110;
		pixels[268*246-1:267*246]=246'b010101001111101011101010101001011111101111111111111111111111111111111111111111111111111111111111111111111111111111111011111101111111111111111111111111111111111111011111111111111101011101011010101101010011010101001011011110111010110101101011010011;
		pixels[269*246-1:268*246]=246'b101010110010010101010101010110111101111111111111111110111110111101111110111111111111111111111111101101111101110111111111111111111111111111101111111111110111011011111111111011110111110110110111010101101110101010110100110101010101101101011110101100;
		pixels[270*246-1:269*246]=246'b010101101101101110101010101101010111111111111111111111101111111111011111111111110111111011111111111111110111111101111111111111111111111011111111111111111111111111111011011110101110101101101100111011011001110000101011101010101011011010110001011011;
		pixels[271*246-1:270*246]=246'b101101010101011011010101010111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111101110111111111110111011111111111111011111111111111011110110101011001101010110001010101101010101010101010111011111101010;
		pixels[272*246-1:271*246]=246'b010101010101101001101010101001011111111111111111101111111111111111111111111111111111011111111111011011011111011111101110110110111111111111111111111111011101111101111111101011011101011011011010110110111011100101010101010101011110111001100100101101;
		pixels[273*246-1:272*246]=246'b101010101010110111010101010111011111111111111011111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111101111111111111111101111110110111111110110110110110111010101100101010010101010101010110101100111011011011010;
		pixels[274*246-1:273*246]=246'b010101010101101100101101010100111111111111111111111111111111111111111111111111011111111111111111111111111111111111111011111111111011010110111011101111111111111111111111110110101101101101101100101101011010101101010101010111101011011100110110110011;
		pixels[275*246-1:274*246]=246'b101101010101111011010010101111011111011101111111111111111111111111111011101111111101110110110111111111111011111011111111011011011111111101111111111101110111111010101101101101111011010101010111110110101101010010101111111001011100101011011010101100;
		pixels[276*246-1:275*246]=246'b110101011010101101101101010010111101111111111111111111111111101111111111111111111111111111111110111111101111111111011111111111110110110111111110111111111110101111111111111110101101110110110010010011010110101001010000101110100111110101101011010111;
		pixels[277*246-1:276*246]=246'b010101010101011010011010101011011111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111101011110111011111111111110110101011110110101101101101101110110101101010101111010101011101001111010110101010;
		pixels[278*246-1:277*246]=246'b101010101011110010110101010110111111111111011111111111111011111110111111111111111111011111111111111111111111011111111111111110111101101101011111011101110101111101011101111110101101011011011011011001101101010100101010110101110010111010101101010101;
		pixels[279*246-1:278*246]=246'b010101010110010110101010101011011111111111111101101110111111111111111111111101101111111011011111101111111111111111111101101111111111111111110111111111111111010111111111010101010110101010101101101110101010101001010101011010101101010101110010111010;
		pixels[280*246-1:279*246]=246'b101010111011101010101101010101111111111111111111111111111111111111111101110111111111111111111011111111111111111111110111111111111111111011111101101110101111111111010101111011111011101101110110110011010101010101011010101101010111011010011101001101;
		pixels[281*246-1:280*246]=246'b010101100100111101011010101110101111110111111111111111111111111111111111111111111011111111111111111111111111111011111111111111101111111110111111111011111101101101111111101110101010011010101010101110101101010100101011010110111010101101100101101010;
		pixels[282*246-1:281*246]=246'b101011011101100001010101101001011111111111111111111111111111101111111111111111111111111111111111111111111011111111111111111111111111111111101110111111110111111011010101010101010101110101101101011001101010101001010110110101100101011011011011011011;
		pixels[283*246-1:282*246]=246'b010101101011011110101010101111111111111110111111111111111111111101110111111111111111111111111111111111111111111111111111111111111110111111111111111110111101011110111110111011101110101010110110101010010101101010101001001010111110100101101101010101;
		pixels[284*246-1:283*246]=246'b011110110101000010110110110010111111011111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111110111101111110111101011010101010010110111010011010111101110110100010110111101001011111110110101101101;
		pixels[285*246-1:284*246]=246'b010010101110111100101101001111011111111111111011011101101101111111011110101111111111111111111111111111111111111111111111111011111111111111111111111111111011011101011101101110111111001100101110110100011001001011010101010011111010101001001011011010;
		pixels[286*246-1:285*246]=246'b101101010100100001011010111001111111111111111111111111111111011111111011111101011011010110111111111111111111110111101110111110111111111111111111111111111110111010110011010101100100111011011000101011110110110100010101101110010101010111110110010111;
		pixels[287*246-1:286*246]=246'b011010101011011110101011001011111111111011011111110111111011110110111111010111110110111111101010110111011101111110111111111111111111111111111111111110111111101111101110111010111011010101100111011101010101001010101010110101101110111010011011101000;
		pixels[288*246-1:287*246]=246'b101011101001000010110101110101111111111111110111111101011111111111101101111010111111101010111111011101110111011111111111101111101101101111111111111111110111110101011011001101001101101010111010100110101010110100000101010110110011001101101100110110;
		pixels[289*246-1:288*246]=246'b010100010110111010101101001011111111111111111110111111101101010101111111101111101010111111011011111111011101110101101010111101110111111010101101101111111110111111110110111011101010101101010101111101010101001011010010101010101110111011010011001000;
		pixels[290*246-1:289*246]=246'b110101111001000101011010110110111101101101011011110111111011111111010101011010010101010101110111010101110111101111011111101011011101010111111011011011011011101010101101010010010101011010101011010010101010110100000101010101011001100010101100010101;


	end
endmodule