module disk200_20(val, pixels);
	input [7:0] val;
	//200*20
	output reg [200*20-1:0] pixels;
	always
	begin
		case(val)		
		1:begin
			pixels[01*200-1:00*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;;
			pixels[02*200-1:01*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[03*200-1:02*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[04*200-1:03*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[05*200-1:04*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[06*200-1:05*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[07*200-1:06*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[08*200-1:07*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[09*200-1:08*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[10*200-1:09*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[11*200-1:10*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[12*200-1:11*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[13*200-1:12*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[14*200-1:13*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[15*200-1:14*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[16*200-1:15*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[17*200-1:16*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[18*200-1:17*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[19*200-1:18*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;
			pixels[20*200-1:19*200]<=200'h0000000000000000000000FFFFFF0000000000000000000000;

		end
		2:begin
			pixels[01*200-1:00*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[02*200-1:01*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[03*200-1:02*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[04*200-1:03*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;			
			pixels[05*200-1:04*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[06*200-1:05*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[07*200-1:06*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[08*200-1:07*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[09*200-1:08*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[10*200-1:09*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[11*200-1:10*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[12*200-1:11*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[13*200-1:12*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[14*200-1:13*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[15*200-1:14*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[16*200-1:15*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[17*200-1:16*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[18*200-1:17*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[19*200-1:18*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;
			pixels[20*200-1:19*200]<=200'h00000000000000000000FFFFFFFFFF00000000000000000000;

		end
		3:begin
			pixels[01*200-1:00*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[02*200-1:01*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[03*200-1:02*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[04*200-1:03*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;			
			pixels[05*200-1:04*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[06*200-1:05*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[07*200-1:06*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[08*200-1:07*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[09*200-1:08*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[10*200-1:09*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[11*200-1:10*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[12*200-1:11*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[13*200-1:12*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[14*200-1:13*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[15*200-1:14*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[16*200-1:15*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[17*200-1:16*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[18*200-1:17*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[19*200-1:18*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;
			pixels[20*200-1:19*200]<=200'h000000000000000000FFFFFFFFFFFFFF000000000000000000;

		end
		4:begin
			pixels[01*200-1:00*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[02*200-1:01*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[03*200-1:02*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[04*200-1:03*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;	
			pixels[05*200-1:04*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[06*200-1:05*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[07*200-1:06*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[08*200-1:07*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[09*200-1:08*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[10*200-1:09*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[11*200-1:10*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[12*200-1:11*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[13*200-1:12*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[14*200-1:13*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[15*200-1:14*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[16*200-1:15*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[17*200-1:16*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[18*200-1:17*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[19*200-1:18*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;
			pixels[20*200-1:19*200]<=200'h0000000000000000FFFFFFFFFFFFFFFFFF0000000000000000;

		end
		5:begin
			pixels[01*200-1:00*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[02*200-1:01*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[03*200-1:02*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[04*200-1:03*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;			
			pixels[05*200-1:04*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[06*200-1:05*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[07*200-1:06*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[08*200-1:07*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[09*200-1:08*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[10*200-1:09*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[11*200-1:10*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[12*200-1:11*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[13*200-1:12*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[14*200-1:13*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[15*200-1:14*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[16*200-1:15*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[17*200-1:16*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[18*200-1:17*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[19*200-1:18*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;
			pixels[20*200-1:19*200]<=200'h00000000000000FFFFFFFFFFFFFFFFFFFFFF00000000000000;

		end
		6:begin
			pixels[01*200-1:00*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[02*200-1:01*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[03*200-1:02*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[04*200-1:03*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;			
			pixels[05*200-1:04*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[06*200-1:05*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[07*200-1:06*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[08*200-1:07*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[09*200-1:08*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[10*200-1:09*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[11*200-1:10*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[12*200-1:11*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[13*200-1:12*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[14*200-1:13*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[15*200-1:14*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[16*200-1:15*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[17*200-1:16*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[18*200-1:17*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[19*200-1:18*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
			pixels[20*200-1:19*200]<=200'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;

		end
		7:begin
			pixels[01*200-1:00*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[02*200-1:01*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[03*200-1:02*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[04*200-1:03*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;			
			pixels[05*200-1:04*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[06*200-1:05*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[07*200-1:06*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[08*200-1:07*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[09*200-1:08*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[10*200-1:09*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[11*200-1:10*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[12*200-1:11*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[13*200-1:12*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[14*200-1:13*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[15*200-1:14*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[16*200-1:15*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[17*200-1:16*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[18*200-1:17*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[19*200-1:18*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
			pixels[20*200-1:19*200]<=200'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;

		end
		8:begin
			pixels[01*200-1:00*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[02*200-1:01*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[03*200-1:02*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[04*200-1:03*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;			
			pixels[05*200-1:04*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[06*200-1:05*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[07*200-1:06*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[08*200-1:07*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[09*200-1:08*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[10*200-1:09*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[11*200-1:10*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[12*200-1:11*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[13*200-1:12*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[14*200-1:13*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[15*200-1:14*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[16*200-1:15*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[17*200-1:16*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[18*200-1:17*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[19*200-1:18*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
			pixels[20*200-1:19*200]<=200'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;

		end
		9:begin
			pixels[01*200-1:00*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[02*200-1:01*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[03*200-1:02*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[04*200-1:03*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;			
			pixels[05*200-1:04*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[06*200-1:05*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[07*200-1:06*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[08*200-1:07*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[09*200-1:08*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[10*200-1:09*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[11*200-1:10*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[12*200-1:11*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[13*200-1:12*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[14*200-1:13*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[15*200-1:14*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[16*200-1:15*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[17*200-1:16*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[18*200-1:17*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[19*200-1:18*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
			pixels[20*200-1:19*200]<=200'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;

		end
		10:begin
			pixels[01*200-1:00*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;			
			pixels[02*200-1:01*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[03*200-1:02*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[04*200-1:03*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;			
			pixels[05*200-1:04*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[06*200-1:05*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[07*200-1:06*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[08*200-1:07*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[09*200-1:08*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[10*200-1:09*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[11*200-1:10*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[12*200-1:11*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[13*200-1:12*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[14*200-1:13*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[15*200-1:14*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[16*200-1:15*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[17*200-1:16*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[18*200-1:17*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[19*200-1:18*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
			pixels[20*200-1:19*200]<=200'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;

		end
		default:begin
			pixels[200*20-1:0]<=4000'b0;
		end
		endcase
		
	end
endmodule