module render(LINE_SEQ, LINE, 
				  DISKa_0, DISKa_1, DISKa_2, DISKa_3, DISKa_4, DISKa_5, DISKa_6, DISKa_7, DISKa_8, DISKa_9,
				  DISKb_0, DISKb_1, DISKb_2, DISKb_3, DISKb_4, DISKb_5, DISKb_6, DISKb_7, DISKb_8, DISKb_9,
				  DISKc_0, DISKc_1, DISKc_2, DISKc_3, DISKc_4, DISKc_5, DISKc_6, DISKc_7, DISKc_8, DISKc_9,
				  TIME_NUM_0, TIME_NUM_1, TIME_NUM_2, TIME_NUM_3,
				  SEL1, SEL2, SEL3,
				  MOVE_NUM_0, MOVE_NUM_1, MOVE_NUM_2, MOVE_NUM_3,

				  BEST_TIME_NUM_0, BEST_TIME_NUM_1, BEST_TIME_NUM_2, BEST_TIME_NUM_3,
				  BEST_MOVE_NUM_0, BEST_MOVE_NUM_1, BEST_MOVE_NUM_2, BEST_MOVE_NUM_3,
				  WON, REC_BREAK_TIME, REC_BREAK_MOVE, M8013
				  );
input [15:0] LINE_SEQ;
output reg [639:0] LINE;
input [7:0] TIME_NUM_0, TIME_NUM_1, TIME_NUM_2, TIME_NUM_3;
input [7:0] MOVE_NUM_0, MOVE_NUM_1, MOVE_NUM_2, MOVE_NUM_3;

input [7:0] BEST_TIME_NUM_0, BEST_TIME_NUM_1, BEST_TIME_NUM_2, BEST_TIME_NUM_3;
input [7:0] BEST_MOVE_NUM_0, BEST_MOVE_NUM_1, BEST_MOVE_NUM_2, BEST_MOVE_NUM_3;

input [7:0] SEL1, SEL2, SEL3;
input [3:0] DISKa_0, DISKa_1, DISKa_2, DISKa_3, DISKa_4, DISKa_5, DISKa_6, DISKa_7, DISKa_8, DISKa_9;
input [3:0] DISKb_0, DISKb_1, DISKb_2, DISKb_3, DISKb_4, DISKb_5, DISKb_6, DISKb_7, DISKb_8, DISKb_9;
input [3:0] DISKc_0, DISKc_1, DISKc_2, DISKc_3, DISKc_4, DISKc_5, DISKc_6, DISKc_7, DISKc_8, DISKc_9;

input WON, REC_BREAK_TIME, REC_BREAK_MOVE, M8013;
//////////////////////////////////////////////////////////////////////////
parameter BEST_B_X = 10, BEST_B_Y = 44;
wire[287:0] BEST_B_PIXMAP;
text12_24 BEST_B_ins(11, BEST_B_PIXMAP);

parameter BEST_E_X = 24, BEST_E_Y = 44;
wire[287:0] BEST_E_PIXMAP;
text12_24 BEST_E_ins(14, BEST_E_PIXMAP);

parameter BEST_S_X = 38, BEST_S_Y = 44;
wire[287:0] BEST_S_PIXMAP;
text12_24 BEST_S_ins(28, BEST_S_PIXMAP);

parameter BEST_T_X = 52, BEST_T_Y = 44;
wire[287:0] BEST_T_PIXMAP;
text12_24 BEST_T_ins(29, BEST_T_PIXMAP);

parameter BEST_DOT_X = 66, BEST_DOT_Y = 44;
wire[287:0] BEST_DOT_PIXMAP;
text12_24 BEST_DOT_ins(36, BEST_DOT_PIXMAP);

//////////////////////////////////////////////////////////////////////////
parameter BEST_TIME_NUM_0_X = 94, BEST_TIME_NUM_0_Y = 44;
wire[287:0] BEST_TIME_NUM_0_PIXMAP;
text12_24 bnum0_ins(BEST_TIME_NUM_0, BEST_TIME_NUM_0_PIXMAP);

parameter BEST_TIME_NUM_1_X = 108, BEST_TIME_NUM_1_Y = 44;
wire[287:0] BEST_TIME_NUM_1_PIXMAP;
text12_24 bnum1_ins(BEST_TIME_NUM_1, BEST_TIME_NUM_1_PIXMAP);

parameter BEST_TIME_NUM_2_X = 136, BEST_TIME_NUM_2_Y = 44;
wire[287:0] BEST_TIME_NUM_2_PIXMAP;
text12_24 bnum2_ins(BEST_TIME_NUM_2, BEST_TIME_NUM_2_PIXMAP);

parameter BEST_TIME_NUM_3_X = 150, BEST_TIME_NUM_3_Y = 44;
wire[287:0] BEST_TIME_NUM_3_PIXMAP;
text12_24 bnum3_ins(BEST_TIME_NUM_3, BEST_TIME_NUM_3_PIXMAP);

//////////////////////////////////////////////////////////////////////////
parameter BEST_MOVE_NUM_0_X = 581, BEST_MOVE_NUM_0_Y = 44;
wire[287:0] BEST_MOVE_NUM_0_PIXMAP;
text12_24 bmove0_ins(BEST_MOVE_NUM_0, BEST_MOVE_NUM_0_PIXMAP);

parameter BEST_MOVE_NUM_1_X = 595, BEST_MOVE_NUM_1_Y = 44;
wire[287:0] BEST_MOVE_NUM_1_PIXMAP;
text12_24 bmove1_ins(BEST_MOVE_NUM_1, BEST_MOVE_NUM_1_PIXMAP);

parameter BEST_MOVE_NUM_2_X = 609, BEST_MOVE_NUM_2_Y = 44;
wire[287:0] BEST_MOVE_NUM_2_PIXMAP;
text12_24 bmove2_ins(BEST_MOVE_NUM_2, BEST_MOVE_NUM_2_PIXMAP);

parameter BEST_MOVE_NUM_3_X = 623, BEST_MOVE_NUM_3_Y = 44;
wire[287:0] BEST_MOVE_NUM_3_PIXMAP;
text12_24 bmove3_ins(BEST_MOVE_NUM_3, BEST_MOVE_NUM_3_PIXMAP);

//////////////////////////////////////////////////////////////////////////
parameter TIME_T_X = 10, TIME_T_Y = 10;
wire[287:0] TIME_T_PIXMAP;
text12_24 NUM_T_ins(29, TIME_T_PIXMAP);

parameter TIME_I_X = 24, TIME_I_Y = 10;
wire[287:0] TIME_I_PIXMAP;
text12_24 NUM_I_ins(18, TIME_I_PIXMAP);

parameter TIME_M_X = 38, TIME_M_Y = 10;
wire[287:0] TIME_M_PIXMAP;
text12_24 NUM_M_ins(22, TIME_M_PIXMAP);

parameter TIME_E_X = 52, TIME_E_Y = 10;
wire[287:0] TIME_E_PIXMAP;
text12_24 NUM_E_ins(14, TIME_E_PIXMAP);

parameter TIME_DOT1_X = 66, TIME_DOT1_Y = 10;
wire[287:0] TIME_DOT1_PIXMAP;
text12_24 NUM_DOT1_ins(36, TIME_DOT1_PIXMAP);


parameter TIME_NUM_0_X = 94, TIME_NUM_0_Y = 10;
wire[287:0] TIME_NUM_0_PIXMAP;
text12_24 num0_ins(TIME_NUM_0, TIME_NUM_0_PIXMAP);

parameter TIME_NUM_1_X = 108, TIME_NUM_1_Y = 10;
wire[287:0] TIME_NUM_1_PIXMAP;
text12_24 num1_ins(TIME_NUM_1, TIME_NUM_1_PIXMAP);

parameter TIME_DOT_X = 122, TIME_DOT_Y = 10;
wire[287:0] TIME_DOT_PIXMAP;
text12_24 NUM_DOT_ins(36, TIME_DOT_PIXMAP);

parameter TIME_NUM_2_X = 136, TIME_NUM_2_Y = 10;
wire[287:0] TIME_NUM_2_PIXMAP;
text12_24 num2_ins(TIME_NUM_2, TIME_NUM_2_PIXMAP);

parameter TIME_NUM_3_X = 150, TIME_NUM_3_Y = 10;
wire[287:0] TIME_NUM_3_PIXMAP;
text12_24 num3_ins(TIME_NUM_3, TIME_NUM_3_PIXMAP);

//////////////////////////////////////////////////////////////////////////
parameter MOVE_M_X = 497, MOVE_M_Y = 10;
wire[287:0] MOVE_M_PIXMAP;
text12_24 MOVE_M_ins(22, MOVE_M_PIXMAP);

parameter MOVE_O_X = 511, MOVE_O_Y = 10;
wire[287:0] MOVE_O_PIXMAP;
text12_24 MOVE_O_ins(24, MOVE_O_PIXMAP);

parameter MOVE_V_X = 525, MOVE_V_Y = 10;
wire[287:0] MOVE_V_PIXMAP;
text12_24 MOVE_V_ins(31, MOVE_V_PIXMAP);

parameter MOVE_E_X = 539, MOVE_E_Y = 10;
wire[287:0] MOVE_E_PIXMAP;
text12_24 MOVE_E_ins(14, MOVE_E_PIXMAP);

parameter MOVE_DOT1_X = 553, MOVE_DOT1_Y = 10;
wire[287:0] MOVE_DOT1_PIXMAP;
text12_24 MOVE_DOT1_ins(36, MOVE_DOT1_PIXMAP);


parameter MOVE_NUM_0_X = 581, MOVE_NUM_0_Y = 10;
wire[287:0] MOVE_NUM_0_PIXMAP;
text12_24 move0_ins(MOVE_NUM_0, MOVE_NUM_0_PIXMAP);

parameter MOVE_NUM_1_X = 595, MOVE_NUM_1_Y = 10;
wire[287:0] MOVE_NUM_1_PIXMAP;
text12_24 move1_ins(MOVE_NUM_1, MOVE_NUM_1_PIXMAP);

parameter MOVE_NUM_2_X = 609, MOVE_NUM_2_Y = 10;
wire[287:0] MOVE_NUM_2_PIXMAP;
text12_24 move2_ins(MOVE_NUM_2, MOVE_NUM_2_PIXMAP);

parameter MOVE_NUM_3_X = 623, MOVE_NUM_3_Y = 10;
wire[287:0] MOVE_NUM_3_PIXMAP;
text12_24 move3_ins(MOVE_NUM_3, MOVE_NUM_3_PIXMAP);

//////////////////////////////////////////////////////////////////////////
parameter SEL1_X = 99, SEL1_Y = 143;
wire[287:0] SEL1_PIXMAP;
text12_24 SEL1_ins(SEL1, SEL1_PIXMAP);

parameter SEL2_X = 314, SEL2_Y = 143;
wire[287:0] SEL2_PIXMAP;
text12_24 SEL2_ins(SEL2, SEL2_PIXMAP);

parameter SEL3_X = 529, SEL3_Y = 143;
wire[287:0] SEL3_PIXMAP;
text12_24 SEL3_ins(SEL3, SEL3_PIXMAP);


//DISKa
//////////////////////////////////////////////////////////////////////////

parameter DISKa_0_X = 5, DISKa_0_Y=430;
wire[4000-1:0] DISKa_0_PIXMAP;
disk200_20 diska_0_ins(DISKa_0, DISKa_0_PIXMAP);

parameter DISKa_1_X = 5, DISKa_1_Y=400;
wire[4000-1:0] DISKa_1_PIXMAP;
disk200_20 diska_1_ins(DISKa_1, DISKa_1_PIXMAP);

parameter DISKa_2_X = 5, DISKa_2_Y=370;
wire[4000-1:0] DISKa_2_PIXMAP;
disk200_20 diska_2_ins(DISKa_2, DISKa_2_PIXMAP);

parameter DISKa_3_X = 5, DISKa_3_Y=340;
wire[4000-1:0] DISKa_3_PIXMAP;
disk200_20 diska_3_ins(DISKa_3, DISKa_3_PIXMAP);

parameter DISKa_4_X = 5, DISKa_4_Y=310;
wire[4000-1:0] DISKa_4_PIXMAP;
disk200_20 diska_4_ins(DISKa_4, DISKa_4_PIXMAP);

parameter DISKa_5_X = 5, DISKa_5_Y=280;
wire[4000-1:0] DISKa_5_PIXMAP;
disk200_20 diska_5_ins(DISKa_5, DISKa_5_PIXMAP);

parameter DISKa_6_X = 5, DISKa_6_Y=250;
wire[4000-1:0] DISKa_6_PIXMAP;
disk200_20 diska_6_ins(DISKa_6, DISKa_6_PIXMAP);

parameter DISKa_7_X = 5, DISKa_7_Y=220;
wire[4000-1:0] DISKa_7_PIXMAP;
disk200_20 diska_7_ins(DISKa_7, DISKa_7_PIXMAP);

parameter DISKa_8_X = 5, DISKa_8_Y=190;
wire[4000-1:0] DISKa_8_PIXMAP;
disk200_20 diska_8_ins(DISKa_8, DISKa_8_PIXMAP);

parameter DISKa_9_X = 5, DISKa_9_Y=160;
wire[4000-1:0] DISKa_9_PIXMAP;
disk200_20 diska_9_ins(DISKa_9, DISKa_9_PIXMAP);
//////////////////////////////////////////////////////////////////////////

//DISKb
//////////////////////////////////////////////////////////////////////////

parameter DISKb_0_X = 220, DISKb_0_Y=430;
wire[4000-1:0] DISKb_0_PIXMAP;
disk200_20 diskb_0_ins(DISKb_0, DISKb_0_PIXMAP);

parameter DISKb_1_X = 220, DISKb_1_Y=400;
wire[4000-1:0] DISKb_1_PIXMAP;
disk200_20 diskb_1_ins(DISKb_1, DISKb_1_PIXMAP);

parameter DISKb_2_X = 220, DISKb_2_Y=370;
wire[4000-1:0] DISKb_2_PIXMAP;
disk200_20 diskb_2_ins(DISKb_2, DISKb_2_PIXMAP);

parameter DISKb_3_X = 220, DISKb_3_Y=340;
wire[4000-1:0] DISKb_3_PIXMAP;
disk200_20 diskb_3_ins(DISKb_3, DISKb_3_PIXMAP);

parameter DISKb_4_X = 220, DISKb_4_Y=310;
wire[4000-1:0] DISKb_4_PIXMAP;
disk200_20 diskb_4_ins(DISKb_4, DISKb_4_PIXMAP);

parameter DISKb_5_X = 220, DISKb_5_Y=280;
wire[4000-1:0] DISKb_5_PIXMAP;
disk200_20 diskb_5_ins(DISKb_5, DISKb_5_PIXMAP);

parameter DISKb_6_X = 220, DISKb_6_Y=250;
wire[4000-1:0] DISKb_6_PIXMAP;
disk200_20 diskb_6_ins(DISKb_6, DISKb_6_PIXMAP);

parameter DISKb_7_X = 220, DISKb_7_Y=220;
wire[4000-1:0] DISKb_7_PIXMAP;
disk200_20 diskb_7_ins(DISKb_7, DISKb_7_PIXMAP);

parameter DISKb_8_X = 220, DISKb_8_Y=190;
wire[4000-1:0] DISKb_8_PIXMAP;
disk200_20 diskb_8_ins(DISKb_8, DISKb_8_PIXMAP);

parameter DISKb_9_X = 220, DISKb_9_Y=160;
wire[4000-1:0] DISKb_9_PIXMAP;
disk200_20 diskb_9_ins(DISKb_9, DISKb_9_PIXMAP);
//////////////////////////////////////////////////////////////////////////

//DISKc
//////////////////////////////////////////////////////////////////////////

parameter DISKc_0_X = 435, DISKc_0_Y=430;
wire[4000-1:0] DISKc_0_PIXMAP;
disk200_20 diskc_0_ins(DISKc_0, DISKc_0_PIXMAP);

parameter DISKc_1_X = 435, DISKc_1_Y=400;
wire[4000-1:0] DISKc_1_PIXMAP;
disk200_20 diskc_1_ins(DISKc_1, DISKc_1_PIXMAP);

parameter DISKc_2_X = 435, DISKc_2_Y=370;
wire[4000-1:0] DISKc_2_PIXMAP;
disk200_20 diskc_2_ins(DISKc_2, DISKc_2_PIXMAP);

parameter DISKc_3_X = 435, DISKc_3_Y=340;
wire[4000-1:0] DISKc_3_PIXMAP;
disk200_20 diskc_3_ins(DISKc_3, DISKc_3_PIXMAP);

parameter DISKc_4_X = 435, DISKc_4_Y=310;
wire[4000-1:0] DISKc_4_PIXMAP;
disk200_20 diskc_4_ins(DISKc_4, DISKc_4_PIXMAP);

parameter DISKc_5_X = 435, DISKc_5_Y=280;
wire[4000-1:0] DISKc_5_PIXMAP;
disk200_20 diskc_5_ins(DISKc_5, DISKc_5_PIXMAP);

parameter DISKc_6_X = 435, DISKc_6_Y=250;
wire[4000-1:0] DISKc_6_PIXMAP;
disk200_20 diskc_6_ins(DISKc_6, DISKc_6_PIXMAP);

parameter DISKc_7_X = 435, DISKc_7_Y=220;
wire[4000-1:0] DISKc_7_PIXMAP;
disk200_20 diskc_7_ins(DISKc_7, DISKc_7_PIXMAP);

parameter DISKc_8_X = 435, DISKc_8_Y=190;
wire[4000-1:0] DISKc_8_PIXMAP;
disk200_20 diskc_8_ins(DISKc_8, DISKc_8_PIXMAP);

parameter DISKc_9_X = 435, DISKc_9_Y=160;
wire[4000-1:0] DISKc_9_PIXMAP;
disk200_20 diskc_9_ins(DISKc_9, DISKc_9_PIXMAP);
//////////////////////////////////////////////////////////////////////////
parameter LAI_0_X = 10, LAI_0_Y = 160;
parameter LAI_1_X = 384, LAI_1_Y = 160;
wire[246*290-1:0] LAI_PIXMAP;
lai246_290 lai_ins(LAI_PIXMAP);

parameter BREAK_RECORD_TIME_X = 188, BREAK_RECORD_TIME_Y = 10;
wire[264*24-1:0] BREAK_RECORD_TIME_PIXMAP;
break_record_time264_24 b_rec_t_ins(BREAK_RECORD_TIME_PIXMAP);

parameter BREAK_RECORD_MOVE_X = 188, BREAK_RECORD_MOVE_Y = 44;
wire[264*24-1:0] BREAK_RECORD_MOVE_PIXMAP;
break_record_move264_24 b_rec_m_ins(BREAK_RECORD_MOVE_PIXMAP);
//////////////////////////////////////////////////////////////////////////
always
begin
	
	
	if(LINE_SEQ==0||LINE_SEQ==479)
	begin		
		LINE<=640'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	end
	else
	begin
		LINE<=640'b0;
		LINE[0]<=1;
		LINE[639]<=1;
	end
	//NUMs
	begin
		if(LINE_SEQ>=TIME_T_Y&&LINE_SEQ<=TIME_T_Y+24)
			render_NUM(LINE_SEQ-TIME_T_Y, LINE[TIME_T_X+12-1:TIME_T_X], TIME_T_PIXMAP);	
		if(LINE_SEQ>=TIME_I_Y&&LINE_SEQ<=TIME_I_Y+24)
			render_NUM(LINE_SEQ-TIME_I_Y, LINE[TIME_I_X+12-1:TIME_I_X], TIME_I_PIXMAP);	
		if(LINE_SEQ>=TIME_M_Y&&LINE_SEQ<=TIME_M_Y+24)
			render_NUM(LINE_SEQ-TIME_M_Y, LINE[TIME_M_X+12-1:TIME_M_X], TIME_M_PIXMAP);	
		if(LINE_SEQ>=TIME_E_Y&&LINE_SEQ<=TIME_E_Y+24)
			render_NUM(LINE_SEQ-TIME_E_Y, LINE[TIME_E_X+12-1:TIME_E_X], TIME_E_PIXMAP);	
		if(LINE_SEQ>=TIME_DOT1_Y&&LINE_SEQ<=TIME_DOT1_Y+24)
			render_NUM(LINE_SEQ-TIME_DOT1_Y, LINE[TIME_DOT1_X+12-1:TIME_DOT1_X], TIME_DOT1_PIXMAP);	
	
		if(LINE_SEQ>=TIME_NUM_0_Y&&LINE_SEQ<=TIME_NUM_0_Y+24)
			render_NUM(LINE_SEQ-TIME_NUM_0_Y, LINE[TIME_NUM_0_X+12-1:TIME_NUM_0_X], TIME_NUM_0_PIXMAP);	
		
		if(LINE_SEQ>=TIME_NUM_1_Y&&LINE_SEQ<=TIME_NUM_1_Y+24)
			render_NUM(LINE_SEQ-TIME_NUM_1_Y, LINE[TIME_NUM_1_X+12-1:TIME_NUM_1_X], TIME_NUM_1_PIXMAP);	
			
		if(LINE_SEQ>=TIME_DOT_Y&&LINE_SEQ<=TIME_DOT_Y+24)
			render_NUM(LINE_SEQ-TIME_DOT_Y, LINE[TIME_DOT_X+12-1:TIME_DOT_X], TIME_DOT_PIXMAP);	
						
		if(LINE_SEQ>=TIME_NUM_2_Y&&LINE_SEQ<=TIME_NUM_2_Y+24)
			render_NUM(LINE_SEQ-TIME_NUM_2_Y, LINE[TIME_NUM_2_X+12-1:TIME_NUM_2_X], TIME_NUM_2_PIXMAP);	
		
		if(LINE_SEQ>=TIME_NUM_3_Y&&LINE_SEQ<=TIME_NUM_3_Y+24)
			render_NUM(LINE_SEQ-TIME_NUM_3_Y, LINE[TIME_NUM_3_X+12-1:TIME_NUM_3_X], TIME_NUM_3_PIXMAP);	
	end
	//MOVEs
	begin
		if(LINE_SEQ>=MOVE_M_Y&&LINE_SEQ<=MOVE_M_Y+24)
			render_NUM(LINE_SEQ-MOVE_M_Y, LINE[MOVE_M_X+12-1:MOVE_M_X], MOVE_M_PIXMAP);	
		if(LINE_SEQ>=MOVE_O_Y&&LINE_SEQ<=MOVE_O_Y+24)
			render_NUM(LINE_SEQ-MOVE_O_Y, LINE[MOVE_O_X+12-1:MOVE_O_X], MOVE_O_PIXMAP);	
		if(LINE_SEQ>=MOVE_V_Y&&LINE_SEQ<=MOVE_V_Y+24)
			render_NUM(LINE_SEQ-MOVE_V_Y, LINE[MOVE_V_X+12-1:MOVE_V_X], MOVE_V_PIXMAP);	
		if(LINE_SEQ>=MOVE_E_Y&&LINE_SEQ<=MOVE_E_Y+24)
			render_NUM(LINE_SEQ-MOVE_E_Y, LINE[MOVE_E_X+12-1:MOVE_E_X], MOVE_E_PIXMAP);	
		if(LINE_SEQ>=MOVE_DOT1_Y&&LINE_SEQ<=MOVE_DOT1_Y+24)
			render_NUM(LINE_SEQ-MOVE_DOT1_Y, LINE[MOVE_DOT1_X+12-1:MOVE_DOT1_X], MOVE_DOT1_PIXMAP);	
	
		if(LINE_SEQ>=MOVE_NUM_0_Y&&LINE_SEQ<=MOVE_NUM_0_Y+24)
			render_NUM(LINE_SEQ-MOVE_NUM_0_Y, LINE[MOVE_NUM_0_X+12-1:MOVE_NUM_0_X], MOVE_NUM_0_PIXMAP);	
		
		if(LINE_SEQ>=MOVE_NUM_1_Y&&LINE_SEQ<=MOVE_NUM_1_Y+24)
			render_NUM(LINE_SEQ-MOVE_NUM_1_Y, LINE[MOVE_NUM_1_X+12-1:MOVE_NUM_1_X], MOVE_NUM_1_PIXMAP);	
			
		if(LINE_SEQ>=MOVE_NUM_2_Y&&LINE_SEQ<=MOVE_NUM_2_Y+24)
			render_NUM(LINE_SEQ-MOVE_NUM_2_Y, LINE[MOVE_NUM_2_X+12-1:MOVE_NUM_2_X], MOVE_NUM_2_PIXMAP);	
		
		if(LINE_SEQ>=MOVE_NUM_3_Y&&LINE_SEQ<=MOVE_NUM_3_Y+24)
			render_NUM(LINE_SEQ-MOVE_NUM_3_Y, LINE[MOVE_NUM_3_X+12-1:MOVE_NUM_3_X], MOVE_NUM_3_PIXMAP);	
	end
	//BEST TIMEs
	begin
		if(LINE_SEQ>=BEST_B_Y&&LINE_SEQ<=BEST_B_Y+24)
			render_NUM(LINE_SEQ-BEST_B_Y, LINE[BEST_B_X+12-1:BEST_B_X], BEST_B_PIXMAP);	
		if(LINE_SEQ>=BEST_E_Y&&LINE_SEQ<=BEST_E_Y+24)
			render_NUM(LINE_SEQ-BEST_E_Y, LINE[BEST_E_X+12-1:BEST_E_X], BEST_E_PIXMAP);	
		if(LINE_SEQ>=BEST_S_Y&&LINE_SEQ<=BEST_S_Y+24)
			render_NUM(LINE_SEQ-BEST_S_Y, LINE[BEST_S_X+12-1:BEST_S_X], BEST_S_PIXMAP);	
		if(LINE_SEQ>=BEST_T_Y&&LINE_SEQ<=BEST_T_Y+24)
			render_NUM(LINE_SEQ-BEST_T_Y, LINE[BEST_T_X+12-1:BEST_T_X], BEST_T_PIXMAP);	
		if(LINE_SEQ>=BEST_DOT_Y&&LINE_SEQ<=BEST_DOT_Y+24)
			render_NUM(LINE_SEQ-BEST_DOT_Y, LINE[BEST_DOT_X+12-1:BEST_DOT_X], BEST_DOT_PIXMAP);	
		
		if(LINE_SEQ>=BEST_DOT_Y&&LINE_SEQ<=BEST_DOT_Y+24)
			render_NUM(LINE_SEQ-BEST_DOT_Y, LINE[BEST_DOT_X+12-1+56:BEST_DOT_X+56], BEST_DOT_PIXMAP);	
			
		if(LINE_SEQ>=BEST_TIME_NUM_0_Y&&LINE_SEQ<=BEST_TIME_NUM_0_Y+24)
			render_NUM(LINE_SEQ-BEST_TIME_NUM_0_Y, LINE[BEST_TIME_NUM_0_X+12-1:BEST_TIME_NUM_0_X], BEST_TIME_NUM_0_PIXMAP);	
		
		if(LINE_SEQ>=BEST_TIME_NUM_1_Y&&LINE_SEQ<=BEST_TIME_NUM_1_Y+24)
			render_NUM(LINE_SEQ-BEST_TIME_NUM_1_Y, LINE[BEST_TIME_NUM_1_X+12-1:BEST_TIME_NUM_1_X], BEST_TIME_NUM_1_PIXMAP);	
						
		if(LINE_SEQ>=BEST_TIME_NUM_2_Y&&LINE_SEQ<=BEST_TIME_NUM_2_Y+24)
			render_NUM(LINE_SEQ-BEST_TIME_NUM_2_Y, LINE[BEST_TIME_NUM_2_X+12-1:BEST_TIME_NUM_2_X], BEST_TIME_NUM_2_PIXMAP);	
		
		if(LINE_SEQ>=BEST_TIME_NUM_3_Y&&LINE_SEQ<=BEST_TIME_NUM_3_Y+24)
			render_NUM(LINE_SEQ-BEST_TIME_NUM_3_Y, LINE[BEST_TIME_NUM_3_X+12-1:BEST_TIME_NUM_3_X], BEST_TIME_NUM_3_PIXMAP);	
	end
	
	//BEST MOVEs	
	begin
		if(LINE_SEQ>=BEST_B_Y&&LINE_SEQ<=BEST_B_Y+24)
			render_NUM(LINE_SEQ-BEST_B_Y, LINE[BEST_B_X+487+12-1:BEST_B_X+487], BEST_B_PIXMAP);	
		if(LINE_SEQ>=BEST_E_Y&&LINE_SEQ<=BEST_E_Y+24)
			render_NUM(LINE_SEQ-BEST_E_Y, LINE[BEST_E_X+487+12-1:BEST_E_X+487], BEST_E_PIXMAP);	
		if(LINE_SEQ>=BEST_S_Y&&LINE_SEQ<=BEST_S_Y+24)
			render_NUM(LINE_SEQ-BEST_S_Y, LINE[BEST_S_X+487+12-1:BEST_S_X+487], BEST_S_PIXMAP);	
		if(LINE_SEQ>=BEST_T_Y&&LINE_SEQ<=BEST_T_Y+24)
			render_NUM(LINE_SEQ-BEST_T_Y, LINE[BEST_T_X+487+12-1:BEST_T_X+487], BEST_T_PIXMAP);	
		if(LINE_SEQ>=BEST_DOT_Y&&LINE_SEQ<=BEST_DOT_Y+24)
			render_NUM(LINE_SEQ-BEST_DOT_Y, LINE[BEST_DOT_X+487+12-1:BEST_DOT_X+487], BEST_DOT_PIXMAP);	
			
		if(LINE_SEQ>=BEST_MOVE_NUM_0_Y&&LINE_SEQ<=BEST_MOVE_NUM_0_Y+24)
			render_NUM(LINE_SEQ-BEST_MOVE_NUM_0_Y, LINE[BEST_MOVE_NUM_0_X+12-1:BEST_MOVE_NUM_0_X], BEST_MOVE_NUM_0_PIXMAP);	
		
		if(LINE_SEQ>=BEST_MOVE_NUM_1_Y&&LINE_SEQ<=BEST_MOVE_NUM_1_Y+24)
			render_NUM(LINE_SEQ-BEST_MOVE_NUM_1_Y, LINE[BEST_MOVE_NUM_1_X+12-1:BEST_MOVE_NUM_1_X], BEST_MOVE_NUM_1_PIXMAP);	
			
		if(LINE_SEQ>=BEST_MOVE_NUM_2_Y&&LINE_SEQ<=BEST_MOVE_NUM_2_Y+24)
			render_NUM(LINE_SEQ-BEST_MOVE_NUM_2_Y, LINE[BEST_MOVE_NUM_2_X+12-1:BEST_MOVE_NUM_2_X], BEST_MOVE_NUM_2_PIXMAP);	
		
		if(LINE_SEQ>=BEST_MOVE_NUM_3_Y&&LINE_SEQ<=BEST_MOVE_NUM_3_Y+24)
			render_NUM(LINE_SEQ-BEST_MOVE_NUM_3_Y, LINE[BEST_MOVE_NUM_3_X+12-1:BEST_MOVE_NUM_3_X], BEST_MOVE_NUM_3_PIXMAP);		
	end

	//SELs
	begin
		if(LINE_SEQ>=SEL1_Y&&LINE_SEQ<=SEL1_Y+24)
			render_NUM(LINE_SEQ-SEL1_Y, LINE[SEL1_X+12-1:SEL1_X], SEL1_PIXMAP);	
			
		if(LINE_SEQ>=SEL2_Y&&LINE_SEQ<=SEL2_Y+24)
			render_NUM(LINE_SEQ-SEL2_Y, LINE[SEL2_X+12-1:SEL2_X], SEL2_PIXMAP);	
			
		if(LINE_SEQ>=SEL3_Y&&LINE_SEQ<=SEL3_Y+24)
			render_NUM(LINE_SEQ-SEL3_Y, LINE[SEL3_X+12-1:SEL3_X], SEL3_PIXMAP);	
	end
	//DISKa	
	begin
		if(LINE_SEQ>=DISKa_0_Y&&LINE_SEQ<=DISKa_0_Y+20)
			render_DISK(LINE_SEQ-DISKa_0_Y, LINE[DISKa_0_X+200-1:DISKa_0_X], DISKa_0_PIXMAP);
		
		if(LINE_SEQ>=DISKa_1_Y&&LINE_SEQ<=DISKa_1_Y+20)
			render_DISK(LINE_SEQ-DISKa_1_Y, LINE[DISKa_1_X+200-1:DISKa_1_X], DISKa_1_PIXMAP);
		
		if(LINE_SEQ>=DISKa_2_Y&&LINE_SEQ<=DISKa_2_Y+20)
			render_DISK(LINE_SEQ-DISKa_2_Y, LINE[DISKa_2_X+200-1:DISKa_2_X], DISKa_2_PIXMAP);
		
		if(LINE_SEQ>=DISKa_3_Y&&LINE_SEQ<=DISKa_3_Y+20)
			render_DISK(LINE_SEQ-DISKa_3_Y, LINE[DISKa_3_X+200-1:DISKa_3_X], DISKa_3_PIXMAP);
		
		if(LINE_SEQ>=DISKa_4_Y&&LINE_SEQ<=DISKa_4_Y+20)
			render_DISK(LINE_SEQ-DISKa_4_Y, LINE[DISKa_4_X+200-1:DISKa_4_X], DISKa_4_PIXMAP);
		
		if(LINE_SEQ>=DISKa_5_Y&&LINE_SEQ<=DISKa_5_Y+20)
			render_DISK(LINE_SEQ-DISKa_5_Y, LINE[DISKa_5_X+200-1:DISKa_5_X], DISKa_5_PIXMAP);
		
		if(LINE_SEQ>=DISKa_6_Y&&LINE_SEQ<=DISKa_6_Y+20)
			render_DISK(LINE_SEQ-DISKa_6_Y, LINE[DISKa_6_X+200-1:DISKa_6_X], DISKa_6_PIXMAP);
		
		if(LINE_SEQ>=DISKa_7_Y&&LINE_SEQ<=DISKa_7_Y+20)
			render_DISK(LINE_SEQ-DISKa_7_Y, LINE[DISKa_7_X+200-1:DISKa_7_X], DISKa_7_PIXMAP);
		
		if(LINE_SEQ>=DISKa_8_Y&&LINE_SEQ<=DISKa_8_Y+20)
			render_DISK(LINE_SEQ-DISKa_8_Y, LINE[DISKa_8_X+200-1:DISKa_8_X], DISKa_8_PIXMAP);
		
		if(LINE_SEQ>=DISKa_9_Y&&LINE_SEQ<=DISKa_9_Y+20)
			render_DISK(LINE_SEQ-DISKa_9_Y, LINE[DISKa_9_X+200-1:DISKa_9_X], DISKa_9_PIXMAP);
	end
	//DISKb	
	begin
		if(LINE_SEQ>=DISKb_0_Y&&LINE_SEQ<=DISKb_0_Y+20)
			render_DISK(LINE_SEQ-DISKb_0_Y, LINE[DISKb_0_X+200-1:DISKb_0_X], DISKb_0_PIXMAP);
		
		if(LINE_SEQ>=DISKb_1_Y&&LINE_SEQ<=DISKb_1_Y+20)
			render_DISK(LINE_SEQ-DISKb_1_Y, LINE[DISKb_1_X+200-1:DISKb_1_X], DISKb_1_PIXMAP);
		
		if(LINE_SEQ>=DISKb_2_Y&&LINE_SEQ<=DISKb_2_Y+20)
			render_DISK(LINE_SEQ-DISKb_2_Y, LINE[DISKb_2_X+200-1:DISKb_2_X], DISKb_2_PIXMAP);
		
		if(LINE_SEQ>=DISKb_3_Y&&LINE_SEQ<=DISKb_3_Y+20)
			render_DISK(LINE_SEQ-DISKb_3_Y, LINE[DISKb_3_X+200-1:DISKb_3_X], DISKb_3_PIXMAP);
		
		if(LINE_SEQ>=DISKb_4_Y&&LINE_SEQ<=DISKb_4_Y+20)
			render_DISK(LINE_SEQ-DISKb_4_Y, LINE[DISKb_4_X+200-1:DISKb_4_X], DISKb_4_PIXMAP);
		
		if(LINE_SEQ>=DISKb_5_Y&&LINE_SEQ<=DISKb_5_Y+20)
			render_DISK(LINE_SEQ-DISKb_5_Y, LINE[DISKb_5_X+200-1:DISKb_5_X], DISKb_5_PIXMAP);
		
		if(LINE_SEQ>=DISKb_6_Y&&LINE_SEQ<=DISKb_6_Y+20)
			render_DISK(LINE_SEQ-DISKb_6_Y, LINE[DISKb_6_X+200-1:DISKb_6_X], DISKb_6_PIXMAP);
		
		if(LINE_SEQ>=DISKb_7_Y&&LINE_SEQ<=DISKb_7_Y+20)
			render_DISK(LINE_SEQ-DISKb_7_Y, LINE[DISKb_7_X+200-1:DISKb_7_X], DISKb_7_PIXMAP);
		
		if(LINE_SEQ>=DISKb_8_Y&&LINE_SEQ<=DISKb_8_Y+20)
			render_DISK(LINE_SEQ-DISKb_8_Y, LINE[DISKb_8_X+200-1:DISKb_8_X], DISKb_8_PIXMAP);
		
		if(LINE_SEQ>=DISKb_9_Y&&LINE_SEQ<=DISKb_9_Y+20)
			render_DISK(LINE_SEQ-DISKb_9_Y, LINE[DISKb_9_X+200-1:DISKb_9_X], DISKb_9_PIXMAP);
	end
	//DISKc	
	begin
		if(LINE_SEQ>=DISKc_0_Y&&LINE_SEQ<=DISKc_0_Y+20)
			render_DISK(LINE_SEQ-DISKc_0_Y, LINE[DISKc_0_X+200-1:DISKc_0_X], DISKc_0_PIXMAP);
		
		if(LINE_SEQ>=DISKc_1_Y&&LINE_SEQ<=DISKc_1_Y+20)
			render_DISK(LINE_SEQ-DISKc_1_Y, LINE[DISKc_1_X+200-1:DISKc_1_X], DISKc_1_PIXMAP);
		
		if(LINE_SEQ>=DISKc_2_Y&&LINE_SEQ<=DISKc_2_Y+20)
			render_DISK(LINE_SEQ-DISKc_2_Y, LINE[DISKc_2_X+200-1:DISKc_2_X], DISKc_2_PIXMAP);
		
		if(LINE_SEQ>=DISKc_3_Y&&LINE_SEQ<=DISKc_3_Y+20)
			render_DISK(LINE_SEQ-DISKc_3_Y, LINE[DISKc_3_X+200-1:DISKc_3_X], DISKc_3_PIXMAP);
		
		if(LINE_SEQ>=DISKc_4_Y&&LINE_SEQ<=DISKc_4_Y+20)
			render_DISK(LINE_SEQ-DISKc_4_Y, LINE[DISKc_4_X+200-1:DISKc_4_X], DISKc_4_PIXMAP);
		
		if(LINE_SEQ>=DISKc_5_Y&&LINE_SEQ<=DISKc_5_Y+20)
			render_DISK(LINE_SEQ-DISKc_5_Y, LINE[DISKc_5_X+200-1:DISKc_5_X], DISKc_5_PIXMAP);
		
		if(LINE_SEQ>=DISKc_6_Y&&LINE_SEQ<=DISKc_6_Y+20)
			render_DISK(LINE_SEQ-DISKc_6_Y, LINE[DISKc_6_X+200-1:DISKc_6_X], DISKc_6_PIXMAP);
		
		if(LINE_SEQ>=DISKc_7_Y&&LINE_SEQ<=DISKc_7_Y+20)
			render_DISK(LINE_SEQ-DISKc_7_Y, LINE[DISKc_7_X+200-1:DISKc_7_X], DISKc_7_PIXMAP);
		
		if(LINE_SEQ>=DISKc_8_Y&&LINE_SEQ<=DISKc_8_Y+20)
			render_DISK(LINE_SEQ-DISKc_8_Y, LINE[DISKc_8_X+200-1:DISKc_8_X], DISKc_8_PIXMAP);
		
		if(LINE_SEQ>=DISKc_9_Y&&LINE_SEQ<=DISKc_9_Y+20)
			render_DISK(LINE_SEQ-DISKc_9_Y, LINE[DISKc_9_X+200-1:DISKc_9_X], DISKc_9_PIXMAP);
	end	
	//WON
	if(WON)
	begin
		if(LINE_SEQ>=LAI_1_Y&&LINE_SEQ<=LAI_1_Y+290&&M8013)
			render_LAI(LINE_SEQ-LAI_1_Y, LINE[LAI_1_X+246-1:LAI_1_X], LAI_PIXMAP);
		if(LINE_SEQ>=LAI_0_Y&&LINE_SEQ<=LAI_0_Y+290&&!M8013)
			render_LAI(LINE_SEQ-LAI_0_Y, LINE[LAI_0_X+246-1:LAI_0_X], LAI_PIXMAP);
		if(M8013&&REC_BREAK_TIME)
		begin
			if(LINE_SEQ>=BREAK_RECORD_TIME_Y&&LINE_SEQ<=BREAK_RECORD_TIME_Y+24)
				render_BREAK_RECORD(LINE_SEQ-BREAK_RECORD_TIME_Y, LINE[BREAK_RECORD_TIME_X+264-1:BREAK_RECORD_TIME_X], BREAK_RECORD_TIME_PIXMAP);
		end
		if(!M8013&&REC_BREAK_MOVE)
		begin
			if(LINE_SEQ>=BREAK_RECORD_MOVE_Y&&LINE_SEQ<=BREAK_RECORD_MOVE_Y+24)
				render_BREAK_RECORD(LINE_SEQ-BREAK_RECORD_MOVE_Y, LINE[BREAK_RECORD_MOVE_X+264-1:BREAK_RECORD_MOVE_X], BREAK_RECORD_MOVE_PIXMAP);
		end
	end
end


task render_DISK;
input [15:0] inY;
output reg [199:0] TARGET;
input [20*200-1:0] PIXMAP;

begin
	case(inY)
				0:	   TARGET=PIXMAP[01*200-1:00*200];
				1:	   TARGET=PIXMAP[02*200-1:01*200];
				2:	   TARGET=PIXMAP[03*200-1:02*200];
				3:	   TARGET=PIXMAP[04*200-1:03*200];
				4:	   TARGET=PIXMAP[05*200-1:04*200];
				5:	   TARGET=PIXMAP[06*200-1:05*200];
				6:	   TARGET=PIXMAP[07*200-1:06*200];
				7:	   TARGET=PIXMAP[08*200-1:07*200];
				8:	   TARGET=PIXMAP[09*200-1:08*200];
				9:	   TARGET=PIXMAP[10*200-1:09*200];
				10:	TARGET=PIXMAP[11*200-1:10*200];
				11:	TARGET=PIXMAP[12*200-1:11*200];
				12:	TARGET=PIXMAP[13*200-1:12*200];
				13:	TARGET=PIXMAP[14*200-1:13*200];
				14:	TARGET=PIXMAP[15*200-1:14*200];
				15:	TARGET=PIXMAP[16*200-1:15*200];
				16:	TARGET=PIXMAP[17*200-1:16*200];
				17:	TARGET=PIXMAP[18*200-1:17*200];
				18:	TARGET=PIXMAP[19*200-1:18*200];
				19:	TARGET=PIXMAP[20*200-1:19*200];
			endcase
end
endtask

task render_NUM;
input [15:0] inY;
output reg [11:0] TARGET;
input [12*24-1:0] PIXMAP;

begin
	case(inY)
				0:	   TARGET=PIXMAP[01*12-1:00*12];
				1:	   TARGET=PIXMAP[02*12-1:01*12];
				2:	   TARGET=PIXMAP[03*12-1:02*12];
				3:	   TARGET=PIXMAP[04*12-1:03*12];
				4:	   TARGET=PIXMAP[05*12-1:04*12];
				5:	   TARGET=PIXMAP[06*12-1:05*12];
				6:	   TARGET=PIXMAP[07*12-1:06*12];
				7:	   TARGET=PIXMAP[08*12-1:07*12];
				8:	   TARGET=PIXMAP[09*12-1:08*12];
				9:	   TARGET=PIXMAP[10*12-1:09*12];
				10:	TARGET=PIXMAP[11*12-1:10*12];
				11:   TARGET=PIXMAP[12*12-1:11*12];
				12:	TARGET=PIXMAP[13*12-1:12*12];
				13:	TARGET=PIXMAP[14*12-1:13*12];
				14:	TARGET=PIXMAP[15*12-1:14*12];
				15:   TARGET=PIXMAP[16*12-1:15*12];
				16:	TARGET=PIXMAP[17*12-1:16*12];
				17:	TARGET=PIXMAP[18*12-1:17*12];
				18:	TARGET=PIXMAP[19*12-1:18*12];
				19:	TARGET=PIXMAP[20*12-1:19*12];
				20:	TARGET=PIXMAP[21*12-1:20*12];
				21:	TARGET=PIXMAP[22*12-1:21*12];
				22:	TARGET=PIXMAP[23*12-1:22*12];
				23:	TARGET=PIXMAP[24*12-1:23*12];
			endcase
end
endtask

task render_LAI;
input [15:0] inY;
output reg [246-1:0] TARGET;
input [246*290-1:0] PIXMAP;

begin
	case(inY)
			0:	   TARGET=PIXMAP[1*246-1:0*246];
			1:	   TARGET=PIXMAP[2*246-1:1*246];
			2:	   TARGET=PIXMAP[3*246-1:2*246];
			3:	   TARGET=PIXMAP[4*246-1:3*246];
			4:	   TARGET=PIXMAP[5*246-1:4*246];
			5:	   TARGET=PIXMAP[6*246-1:5*246];
			6:	   TARGET=PIXMAP[7*246-1:6*246];
			7:	   TARGET=PIXMAP[8*246-1:7*246];
			8:	   TARGET=PIXMAP[9*246-1:8*246];
			9:	   TARGET=PIXMAP[10*246-1:9*246];
			10:	   TARGET=PIXMAP[11*246-1:10*246];
			11:	   TARGET=PIXMAP[12*246-1:11*246];
			12:	   TARGET=PIXMAP[13*246-1:12*246];
			13:	   TARGET=PIXMAP[14*246-1:13*246];
			14:	   TARGET=PIXMAP[15*246-1:14*246];
			15:	   TARGET=PIXMAP[16*246-1:15*246];
			16:	   TARGET=PIXMAP[17*246-1:16*246];
			17:	   TARGET=PIXMAP[18*246-1:17*246];
			18:	   TARGET=PIXMAP[19*246-1:18*246];
			19:	   TARGET=PIXMAP[20*246-1:19*246];
			20:	   TARGET=PIXMAP[21*246-1:20*246];
			21:	   TARGET=PIXMAP[22*246-1:21*246];
			22:	   TARGET=PIXMAP[23*246-1:22*246];
			23:	   TARGET=PIXMAP[24*246-1:23*246];
			24:	   TARGET=PIXMAP[25*246-1:24*246];
			25:	   TARGET=PIXMAP[26*246-1:25*246];
			26:	   TARGET=PIXMAP[27*246-1:26*246];
			27:	   TARGET=PIXMAP[28*246-1:27*246];
			28:	   TARGET=PIXMAP[29*246-1:28*246];
			29:	   TARGET=PIXMAP[30*246-1:29*246];
			30:	   TARGET=PIXMAP[31*246-1:30*246];
			31:	   TARGET=PIXMAP[32*246-1:31*246];
			32:	   TARGET=PIXMAP[33*246-1:32*246];
			33:	   TARGET=PIXMAP[34*246-1:33*246];
			34:	   TARGET=PIXMAP[35*246-1:34*246];
			35:	   TARGET=PIXMAP[36*246-1:35*246];
			36:	   TARGET=PIXMAP[37*246-1:36*246];
			37:	   TARGET=PIXMAP[38*246-1:37*246];
			38:	   TARGET=PIXMAP[39*246-1:38*246];
			39:	   TARGET=PIXMAP[40*246-1:39*246];
			40:	   TARGET=PIXMAP[41*246-1:40*246];
			41:	   TARGET=PIXMAP[42*246-1:41*246];
			42:	   TARGET=PIXMAP[43*246-1:42*246];
			43:	   TARGET=PIXMAP[44*246-1:43*246];
			44:	   TARGET=PIXMAP[45*246-1:44*246];
			45:	   TARGET=PIXMAP[46*246-1:45*246];
			46:	   TARGET=PIXMAP[47*246-1:46*246];
			47:	   TARGET=PIXMAP[48*246-1:47*246];
			48:	   TARGET=PIXMAP[49*246-1:48*246];
			49:	   TARGET=PIXMAP[50*246-1:49*246];
			50:	   TARGET=PIXMAP[51*246-1:50*246];
			51:	   TARGET=PIXMAP[52*246-1:51*246];
			52:	   TARGET=PIXMAP[53*246-1:52*246];
			53:	   TARGET=PIXMAP[54*246-1:53*246];
			54:	   TARGET=PIXMAP[55*246-1:54*246];
			55:	   TARGET=PIXMAP[56*246-1:55*246];
			56:	   TARGET=PIXMAP[57*246-1:56*246];
			57:	   TARGET=PIXMAP[58*246-1:57*246];
			58:	   TARGET=PIXMAP[59*246-1:58*246];
			59:	   TARGET=PIXMAP[60*246-1:59*246];
			60:	   TARGET=PIXMAP[61*246-1:60*246];
			61:	   TARGET=PIXMAP[62*246-1:61*246];
			62:	   TARGET=PIXMAP[63*246-1:62*246];
			63:	   TARGET=PIXMAP[64*246-1:63*246];
			64:	   TARGET=PIXMAP[65*246-1:64*246];
			65:	   TARGET=PIXMAP[66*246-1:65*246];
			66:	   TARGET=PIXMAP[67*246-1:66*246];
			67:	   TARGET=PIXMAP[68*246-1:67*246];
			68:	   TARGET=PIXMAP[69*246-1:68*246];
			69:	   TARGET=PIXMAP[70*246-1:69*246];
			70:	   TARGET=PIXMAP[71*246-1:70*246];
			71:	   TARGET=PIXMAP[72*246-1:71*246];
			72:	   TARGET=PIXMAP[73*246-1:72*246];
			73:	   TARGET=PIXMAP[74*246-1:73*246];
			74:	   TARGET=PIXMAP[75*246-1:74*246];
			75:	   TARGET=PIXMAP[76*246-1:75*246];
			76:	   TARGET=PIXMAP[77*246-1:76*246];
			77:	   TARGET=PIXMAP[78*246-1:77*246];
			78:	   TARGET=PIXMAP[79*246-1:78*246];
			79:	   TARGET=PIXMAP[80*246-1:79*246];
			80:	   TARGET=PIXMAP[81*246-1:80*246];
			81:	   TARGET=PIXMAP[82*246-1:81*246];
			82:	   TARGET=PIXMAP[83*246-1:82*246];
			83:	   TARGET=PIXMAP[84*246-1:83*246];
			84:	   TARGET=PIXMAP[85*246-1:84*246];
			85:	   TARGET=PIXMAP[86*246-1:85*246];
			86:	   TARGET=PIXMAP[87*246-1:86*246];
			87:	   TARGET=PIXMAP[88*246-1:87*246];
			88:	   TARGET=PIXMAP[89*246-1:88*246];
			89:	   TARGET=PIXMAP[90*246-1:89*246];
			90:	   TARGET=PIXMAP[91*246-1:90*246];
			91:	   TARGET=PIXMAP[92*246-1:91*246];
			92:	   TARGET=PIXMAP[93*246-1:92*246];
			93:	   TARGET=PIXMAP[94*246-1:93*246];
			94:	   TARGET=PIXMAP[95*246-1:94*246];
			95:	   TARGET=PIXMAP[96*246-1:95*246];
			96:	   TARGET=PIXMAP[97*246-1:96*246];
			97:	   TARGET=PIXMAP[98*246-1:97*246];
			98:	   TARGET=PIXMAP[99*246-1:98*246];
			99:	   TARGET=PIXMAP[100*246-1:99*246];
			100:	   TARGET=PIXMAP[101*246-1:100*246];
			101:	   TARGET=PIXMAP[102*246-1:101*246];
			102:	   TARGET=PIXMAP[103*246-1:102*246];
			103:	   TARGET=PIXMAP[104*246-1:103*246];
			104:	   TARGET=PIXMAP[105*246-1:104*246];
			105:	   TARGET=PIXMAP[106*246-1:105*246];
			106:	   TARGET=PIXMAP[107*246-1:106*246];
			107:	   TARGET=PIXMAP[108*246-1:107*246];
			108:	   TARGET=PIXMAP[109*246-1:108*246];
			109:	   TARGET=PIXMAP[110*246-1:109*246];
			110:	   TARGET=PIXMAP[111*246-1:110*246];
			111:	   TARGET=PIXMAP[112*246-1:111*246];
			112:	   TARGET=PIXMAP[113*246-1:112*246];
			113:	   TARGET=PIXMAP[114*246-1:113*246];
			114:	   TARGET=PIXMAP[115*246-1:114*246];
			115:	   TARGET=PIXMAP[116*246-1:115*246];
			116:	   TARGET=PIXMAP[117*246-1:116*246];
			117:	   TARGET=PIXMAP[118*246-1:117*246];
			118:	   TARGET=PIXMAP[119*246-1:118*246];
			119:	   TARGET=PIXMAP[120*246-1:119*246];
			120:	   TARGET=PIXMAP[121*246-1:120*246];
			121:	   TARGET=PIXMAP[122*246-1:121*246];
			122:	   TARGET=PIXMAP[123*246-1:122*246];
			123:	   TARGET=PIXMAP[124*246-1:123*246];
			124:	   TARGET=PIXMAP[125*246-1:124*246];
			125:	   TARGET=PIXMAP[126*246-1:125*246];
			126:	   TARGET=PIXMAP[127*246-1:126*246];
			127:	   TARGET=PIXMAP[128*246-1:127*246];
			128:	   TARGET=PIXMAP[129*246-1:128*246];
			129:	   TARGET=PIXMAP[130*246-1:129*246];
			130:	   TARGET=PIXMAP[131*246-1:130*246];
			131:	   TARGET=PIXMAP[132*246-1:131*246];
			132:	   TARGET=PIXMAP[133*246-1:132*246];
			133:	   TARGET=PIXMAP[134*246-1:133*246];
			134:	   TARGET=PIXMAP[135*246-1:134*246];
			135:	   TARGET=PIXMAP[136*246-1:135*246];
			136:	   TARGET=PIXMAP[137*246-1:136*246];
			137:	   TARGET=PIXMAP[138*246-1:137*246];
			138:	   TARGET=PIXMAP[139*246-1:138*246];
			139:	   TARGET=PIXMAP[140*246-1:139*246];
			140:	   TARGET=PIXMAP[141*246-1:140*246];
			141:	   TARGET=PIXMAP[142*246-1:141*246];
			142:	   TARGET=PIXMAP[143*246-1:142*246];
			143:	   TARGET=PIXMAP[144*246-1:143*246];
			144:	   TARGET=PIXMAP[145*246-1:144*246];
			145:	   TARGET=PIXMAP[146*246-1:145*246];
			146:	   TARGET=PIXMAP[147*246-1:146*246];
			147:	   TARGET=PIXMAP[148*246-1:147*246];
			148:	   TARGET=PIXMAP[149*246-1:148*246];
			149:	   TARGET=PIXMAP[150*246-1:149*246];
			150:	   TARGET=PIXMAP[151*246-1:150*246];
			151:	   TARGET=PIXMAP[152*246-1:151*246];
			152:	   TARGET=PIXMAP[153*246-1:152*246];
			153:	   TARGET=PIXMAP[154*246-1:153*246];
			154:	   TARGET=PIXMAP[155*246-1:154*246];
			155:	   TARGET=PIXMAP[156*246-1:155*246];
			156:	   TARGET=PIXMAP[157*246-1:156*246];
			157:	   TARGET=PIXMAP[158*246-1:157*246];
			158:	   TARGET=PIXMAP[159*246-1:158*246];
			159:	   TARGET=PIXMAP[160*246-1:159*246];
			160:	   TARGET=PIXMAP[161*246-1:160*246];
			161:	   TARGET=PIXMAP[162*246-1:161*246];
			162:	   TARGET=PIXMAP[163*246-1:162*246];
			163:	   TARGET=PIXMAP[164*246-1:163*246];
			164:	   TARGET=PIXMAP[165*246-1:164*246];
			165:	   TARGET=PIXMAP[166*246-1:165*246];
			166:	   TARGET=PIXMAP[167*246-1:166*246];
			167:	   TARGET=PIXMAP[168*246-1:167*246];
			168:	   TARGET=PIXMAP[169*246-1:168*246];
			169:	   TARGET=PIXMAP[170*246-1:169*246];
			170:	   TARGET=PIXMAP[171*246-1:170*246];
			171:	   TARGET=PIXMAP[172*246-1:171*246];
			172:	   TARGET=PIXMAP[173*246-1:172*246];
			173:	   TARGET=PIXMAP[174*246-1:173*246];
			174:	   TARGET=PIXMAP[175*246-1:174*246];
			175:	   TARGET=PIXMAP[176*246-1:175*246];
			176:	   TARGET=PIXMAP[177*246-1:176*246];
			177:	   TARGET=PIXMAP[178*246-1:177*246];
			178:	   TARGET=PIXMAP[179*246-1:178*246];
			179:	   TARGET=PIXMAP[180*246-1:179*246];
			180:	   TARGET=PIXMAP[181*246-1:180*246];
			181:	   TARGET=PIXMAP[182*246-1:181*246];
			182:	   TARGET=PIXMAP[183*246-1:182*246];
			183:	   TARGET=PIXMAP[184*246-1:183*246];
			184:	   TARGET=PIXMAP[185*246-1:184*246];
			185:	   TARGET=PIXMAP[186*246-1:185*246];
			186:	   TARGET=PIXMAP[187*246-1:186*246];
			187:	   TARGET=PIXMAP[188*246-1:187*246];
			188:	   TARGET=PIXMAP[189*246-1:188*246];
			189:	   TARGET=PIXMAP[190*246-1:189*246];
			190:	   TARGET=PIXMAP[191*246-1:190*246];
			191:	   TARGET=PIXMAP[192*246-1:191*246];
			192:	   TARGET=PIXMAP[193*246-1:192*246];
			193:	   TARGET=PIXMAP[194*246-1:193*246];
			194:	   TARGET=PIXMAP[195*246-1:194*246];
			195:	   TARGET=PIXMAP[196*246-1:195*246];
			196:	   TARGET=PIXMAP[197*246-1:196*246];
			197:	   TARGET=PIXMAP[198*246-1:197*246];
			198:	   TARGET=PIXMAP[199*246-1:198*246];
			199:	   TARGET=PIXMAP[200*246-1:199*246];
			200:	   TARGET=PIXMAP[201*246-1:200*246];
			201:	   TARGET=PIXMAP[202*246-1:201*246];
			202:	   TARGET=PIXMAP[203*246-1:202*246];
			203:	   TARGET=PIXMAP[204*246-1:203*246];
			204:	   TARGET=PIXMAP[205*246-1:204*246];
			205:	   TARGET=PIXMAP[206*246-1:205*246];
			206:	   TARGET=PIXMAP[207*246-1:206*246];
			207:	   TARGET=PIXMAP[208*246-1:207*246];
			208:	   TARGET=PIXMAP[209*246-1:208*246];
			209:	   TARGET=PIXMAP[210*246-1:209*246];
			210:	   TARGET=PIXMAP[211*246-1:210*246];
			211:	   TARGET=PIXMAP[212*246-1:211*246];
			212:	   TARGET=PIXMAP[213*246-1:212*246];
			213:	   TARGET=PIXMAP[214*246-1:213*246];
			214:	   TARGET=PIXMAP[215*246-1:214*246];
			215:	   TARGET=PIXMAP[216*246-1:215*246];
			216:	   TARGET=PIXMAP[217*246-1:216*246];
			217:	   TARGET=PIXMAP[218*246-1:217*246];
			218:	   TARGET=PIXMAP[219*246-1:218*246];
			219:	   TARGET=PIXMAP[220*246-1:219*246];
			220:	   TARGET=PIXMAP[221*246-1:220*246];
			221:	   TARGET=PIXMAP[222*246-1:221*246];
			222:	   TARGET=PIXMAP[223*246-1:222*246];
			223:	   TARGET=PIXMAP[224*246-1:223*246];
			224:	   TARGET=PIXMAP[225*246-1:224*246];
			225:	   TARGET=PIXMAP[226*246-1:225*246];
			226:	   TARGET=PIXMAP[227*246-1:226*246];
			227:	   TARGET=PIXMAP[228*246-1:227*246];
			228:	   TARGET=PIXMAP[229*246-1:228*246];
			229:	   TARGET=PIXMAP[230*246-1:229*246];
			230:	   TARGET=PIXMAP[231*246-1:230*246];
			231:	   TARGET=PIXMAP[232*246-1:231*246];
			232:	   TARGET=PIXMAP[233*246-1:232*246];
			233:	   TARGET=PIXMAP[234*246-1:233*246];
			234:	   TARGET=PIXMAP[235*246-1:234*246];
			235:	   TARGET=PIXMAP[236*246-1:235*246];
			236:	   TARGET=PIXMAP[237*246-1:236*246];
			237:	   TARGET=PIXMAP[238*246-1:237*246];
			238:	   TARGET=PIXMAP[239*246-1:238*246];
			239:	   TARGET=PIXMAP[240*246-1:239*246];
			240:	   TARGET=PIXMAP[241*246-1:240*246];
			241:	   TARGET=PIXMAP[242*246-1:241*246];
			242:	   TARGET=PIXMAP[243*246-1:242*246];
			243:	   TARGET=PIXMAP[244*246-1:243*246];
			244:	   TARGET=PIXMAP[245*246-1:244*246];
			245:	   TARGET=PIXMAP[246*246-1:245*246];
			246:	   TARGET=PIXMAP[247*246-1:246*246];
			247:	   TARGET=PIXMAP[248*246-1:247*246];
			248:	   TARGET=PIXMAP[249*246-1:248*246];
			249:	   TARGET=PIXMAP[250*246-1:249*246];
			250:	   TARGET=PIXMAP[251*246-1:250*246];
			251:	   TARGET=PIXMAP[252*246-1:251*246];
			252:	   TARGET=PIXMAP[253*246-1:252*246];
			253:	   TARGET=PIXMAP[254*246-1:253*246];
			254:	   TARGET=PIXMAP[255*246-1:254*246];
			255:	   TARGET=PIXMAP[256*246-1:255*246];
			256:	   TARGET=PIXMAP[257*246-1:256*246];
			257:	   TARGET=PIXMAP[258*246-1:257*246];
			258:	   TARGET=PIXMAP[259*246-1:258*246];
			259:	   TARGET=PIXMAP[260*246-1:259*246];
			260:	   TARGET=PIXMAP[261*246-1:260*246];
			261:	   TARGET=PIXMAP[262*246-1:261*246];
			262:	   TARGET=PIXMAP[263*246-1:262*246];
			263:	   TARGET=PIXMAP[264*246-1:263*246];
			264:	   TARGET=PIXMAP[265*246-1:264*246];
			265:	   TARGET=PIXMAP[266*246-1:265*246];
			266:	   TARGET=PIXMAP[267*246-1:266*246];
			267:	   TARGET=PIXMAP[268*246-1:267*246];
			268:	   TARGET=PIXMAP[269*246-1:268*246];
			269:	   TARGET=PIXMAP[270*246-1:269*246];
			270:	   TARGET=PIXMAP[271*246-1:270*246];
			271:	   TARGET=PIXMAP[272*246-1:271*246];
			272:	   TARGET=PIXMAP[273*246-1:272*246];
			273:	   TARGET=PIXMAP[274*246-1:273*246];
			274:	   TARGET=PIXMAP[275*246-1:274*246];
			275:	   TARGET=PIXMAP[276*246-1:275*246];
			276:	   TARGET=PIXMAP[277*246-1:276*246];
			277:	   TARGET=PIXMAP[278*246-1:277*246];
			278:	   TARGET=PIXMAP[279*246-1:278*246];
			279:	   TARGET=PIXMAP[280*246-1:279*246];
			280:	   TARGET=PIXMAP[281*246-1:280*246];
			281:	   TARGET=PIXMAP[282*246-1:281*246];
			282:	   TARGET=PIXMAP[283*246-1:282*246];
			283:	   TARGET=PIXMAP[284*246-1:283*246];
			284:	   TARGET=PIXMAP[285*246-1:284*246];
			285:	   TARGET=PIXMAP[286*246-1:285*246];
			286:	   TARGET=PIXMAP[287*246-1:286*246];
			287:	   TARGET=PIXMAP[288*246-1:287*246];
			288:	   TARGET=PIXMAP[289*246-1:288*246];
			289:	   TARGET=PIXMAP[290*246-1:289*246];
		endcase
end
endtask

task render_BREAK_RECORD;
input [15:0] inY;
output reg [264-1:0] TARGET;
input [264*24-1:0] PIXMAP;

begin
	case(inY)
		0:	      TARGET=PIXMAP[1*264-1:0*264];
		1:	      TARGET=PIXMAP[2*264-1:1*264];
		2:	      TARGET=PIXMAP[3*264-1:2*264];
		3:	      TARGET=PIXMAP[4*264-1:3*264];
		4:	      TARGET=PIXMAP[5*264-1:4*264];
		5:	      TARGET=PIXMAP[6*264-1:5*264];
		6:	      TARGET=PIXMAP[7*264-1:6*264];
		7:	      TARGET=PIXMAP[8*264-1:7*264];
		8:	      TARGET=PIXMAP[9*264-1:8*264];
		9:	      TARGET=PIXMAP[10*264-1:9*264];
		10:	   TARGET=PIXMAP[11*264-1:10*264];
		11:	   TARGET=PIXMAP[12*264-1:11*264];
		12:	   TARGET=PIXMAP[13*264-1:12*264];
		13:	   TARGET=PIXMAP[14*264-1:13*264];
		14:	   TARGET=PIXMAP[15*264-1:14*264];
		15:	   TARGET=PIXMAP[16*264-1:15*264];
		16:	   TARGET=PIXMAP[17*264-1:16*264];
		17:	   TARGET=PIXMAP[18*264-1:17*264];
		18:	   TARGET=PIXMAP[19*264-1:18*264];
		19:	   TARGET=PIXMAP[20*264-1:19*264];
		20:	   TARGET=PIXMAP[21*264-1:20*264];
		21:	   TARGET=PIXMAP[22*264-1:21*264];
		22:	   TARGET=PIXMAP[23*264-1:22*264];
		23:	   TARGET=PIXMAP[24*264-1:23*264];
	endcase
end
endtask

endmodule

