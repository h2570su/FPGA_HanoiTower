module text12_24(val, pixels);
	input [7:0] val;
	//12*24
	output reg [12*24-1:0] pixels;
	always
	begin
		case(val)
		0:begin
			pixels[01*12-1:00*12]<=12'b111111111111;			
			pixels[02*12-1:01*12]<=12'b111111111111;
			pixels[03*12-1:02*12]<=12'b111111111111;
			pixels[04*12-1:03*12]<=12'b111111111111;			
			pixels[05*12-1:04*12]<=12'b111000000111;
			pixels[06*12-1:05*12]<=12'b111000000111;
			pixels[07*12-1:06*12]<=12'b111000000111;
			pixels[08*12-1:07*12]<=12'b111000000111;
			pixels[09*12-1:08*12]<=12'b111000000111;
			pixels[10*12-1:09*12]<=12'b111000000111;
			pixels[11*12-1:10*12]<=12'b111000000111;
			pixels[12*12-1:11*12]<=12'b111000000111;
			pixels[13*12-1:12*12]<=12'b111000000111;
			pixels[14*12-1:13*12]<=12'b111000000111;
			pixels[15*12-1:14*12]<=12'b111000000111;
			pixels[16*12-1:15*12]<=12'b111000000111;
			pixels[17*12-1:16*12]<=12'b111000000111;
			pixels[18*12-1:17*12]<=12'b111000000111;
			pixels[19*12-1:18*12]<=12'b111000000111;
			pixels[20*12-1:19*12]<=12'b111000000111;
			pixels[21*12-1:20*12]<=12'b111111111111;
			pixels[22*12-1:21*12]<=12'b111111111111;
			pixels[23*12-1:22*12]<=12'b111111111111;
			pixels[24*12-1:23*12]<=12'b111111111111;
		end
		1:begin
			pixels[01*12-1:00*12]<=12'b111000000000;
			pixels[02*12-1:01*12]<=12'b111000000000;
			pixels[03*12-1:02*12]<=12'b111000000000;
			pixels[04*12-1:03*12]<=12'b111000000000;
			pixels[05*12-1:04*12]<=12'b111000000000;
			pixels[06*12-1:05*12]<=12'b111000000000;
			pixels[07*12-1:06*12]<=12'b111000000000;
			pixels[08*12-1:07*12]<=12'b111000000000;
			pixels[09*12-1:08*12]<=12'b111000000000;
			pixels[10*12-1:09*12]<=12'b111000000000;
			pixels[11*12-1:10*12]<=12'b111000000000;
			pixels[12*12-1:11*12]<=12'b111000000000;
			pixels[13*12-1:12*12]<=12'b111000000000;
			pixels[14*12-1:13*12]<=12'b111000000000;
			pixels[15*12-1:14*12]<=12'b111000000000;
			pixels[16*12-1:15*12]<=12'b111000000000;
			pixels[17*12-1:16*12]<=12'b111000000000;
			pixels[18*12-1:17*12]<=12'b111000000000;
			pixels[19*12-1:18*12]<=12'b111000000000;
			pixels[20*12-1:19*12]<=12'b111000000000;
			pixels[21*12-1:20*12]<=12'b111000000000;
			pixels[22*12-1:21*12]<=12'b111000000000;
			pixels[23*12-1:22*12]<=12'b111000000000;
			pixels[24*12-1:23*12]<=12'b111000000000;
		end
		2:begin
			pixels[01*12-1:00*12]<=12'b111111111111;
			pixels[02*12-1:01*12]<=12'b111111111111;
			pixels[03*12-1:02*12]<=12'b111111111111;
			pixels[04*12-1:03*12]<=12'b111111111111;			
			pixels[05*12-1:04*12]<=12'b111000000000;
			pixels[06*12-1:05*12]<=12'b111000000000;
			pixels[07*12-1:06*12]<=12'b111000000000;
			pixels[08*12-1:07*12]<=12'b111000000000;
			pixels[09*12-1:08*12]<=12'b111000000000;
			pixels[10*12-1:09*12]<=12'b111000000000;
			pixels[11*12-1:10*12]<=12'b111000000000;
			pixels[12*12-1:11*12]<=12'b111111111111;
			pixels[13*12-1:12*12]<=12'b111111111111;
			pixels[14*12-1:13*12]<=12'b000000000111;
			pixels[15*12-1:14*12]<=12'b000000000111;
			pixels[16*12-1:15*12]<=12'b000000000111;
			pixels[17*12-1:16*12]<=12'b000000000111;
			pixels[18*12-1:17*12]<=12'b000000000111;
			pixels[19*12-1:18*12]<=12'b000000000111;
			pixels[20*12-1:19*12]<=12'b000000000111;
			pixels[21*12-1:20*12]<=12'b111111111111;
			pixels[22*12-1:21*12]<=12'b111111111111;
			pixels[23*12-1:22*12]<=12'b111111111111;
			pixels[24*12-1:23*12]<=12'b111111111111;
		end
		3:begin
			pixels[01*12-1:00*12]<=12'b111111111111;
			pixels[02*12-1:01*12]<=12'b111111111111;
			pixels[03*12-1:02*12]<=12'b111111111111;
			pixels[04*12-1:03*12]<=12'b111111111111;			
			pixels[05*12-1:04*12]<=12'b111000000000;
			pixels[06*12-1:05*12]<=12'b111000000000;
			pixels[07*12-1:06*12]<=12'b111000000000;
			pixels[08*12-1:07*12]<=12'b111000000000;
			pixels[09*12-1:08*12]<=12'b111000000000;
			pixels[10*12-1:09*12]<=12'b111000000000;
			pixels[11*12-1:10*12]<=12'b111000000000;
			pixels[12*12-1:11*12]<=12'b111111111111;
			pixels[13*12-1:12*12]<=12'b111111111111;
			pixels[14*12-1:13*12]<=12'b111000000000;
			pixels[15*12-1:14*12]<=12'b111000000000;
			pixels[16*12-1:15*12]<=12'b111000000000;
			pixels[17*12-1:16*12]<=12'b111000000000;
			pixels[18*12-1:17*12]<=12'b111000000000;
			pixels[19*12-1:18*12]<=12'b111000000000;
			pixels[20*12-1:19*12]<=12'b111000000000;
			pixels[21*12-1:20*12]<=12'b111111111111;
			pixels[22*12-1:21*12]<=12'b111111111111;
			pixels[23*12-1:22*12]<=12'b111111111111;
			pixels[24*12-1:23*12]<=12'b111111111111;
		end
		4:begin
			pixels[01*12-1:00*12]<=12'b111000000111;
			pixels[02*12-1:01*12]<=12'b111000000111;
			pixels[03*12-1:02*12]<=12'b111000000111;
			pixels[04*12-1:03*12]<=12'b111000000111;	
			pixels[05*12-1:04*12]<=12'b111000000111;
			pixels[06*12-1:05*12]<=12'b111000000111;
			pixels[07*12-1:06*12]<=12'b111000000111;
			pixels[08*12-1:07*12]<=12'b111000000111;
			pixels[09*12-1:08*12]<=12'b111000000111;
			pixels[10*12-1:09*12]<=12'b111000000111;
			pixels[11*12-1:10*12]<=12'b111000000111;
			pixels[12*12-1:11*12]<=12'b111111111111;
			pixels[13*12-1:12*12]<=12'b111111111111;
			pixels[14*12-1:13*12]<=12'b111000000000;
			pixels[15*12-1:14*12]<=12'b111000000000;
			pixels[16*12-1:15*12]<=12'b111000000000;
			pixels[17*12-1:16*12]<=12'b111000000000;
			pixels[18*12-1:17*12]<=12'b111000000000;
			pixels[19*12-1:18*12]<=12'b111000000000;
			pixels[20*12-1:19*12]<=12'b111000000000;
			pixels[21*12-1:20*12]<=12'b111000000000;
			pixels[22*12-1:21*12]<=12'b111000000000;
			pixels[23*12-1:22*12]<=12'b111000000000;
			pixels[24*12-1:23*12]<=12'b111000000000;
		end
		5:begin
			pixels[01*12-1:00*12]<=12'b111111111111;
			pixels[02*12-1:01*12]<=12'b111111111111;
			pixels[03*12-1:02*12]<=12'b111111111111;
			pixels[04*12-1:03*12]<=12'b111111111111;			
			pixels[05*12-1:04*12]<=12'b000000000111;
			pixels[06*12-1:05*12]<=12'b000000000111;
			pixels[07*12-1:06*12]<=12'b000000000111;
			pixels[08*12-1:07*12]<=12'b000000000111;
			pixels[09*12-1:08*12]<=12'b000000000111;
			pixels[10*12-1:09*12]<=12'b000000000111;
			pixels[11*12-1:10*12]<=12'b000000000111;
			pixels[12*12-1:11*12]<=12'b111111111111;
			pixels[13*12-1:12*12]<=12'b111111111111;
			pixels[14*12-1:13*12]<=12'b111000000000;
			pixels[15*12-1:14*12]<=12'b111000000000;
			pixels[16*12-1:15*12]<=12'b111000000000;
			pixels[17*12-1:16*12]<=12'b111000000000;
			pixels[18*12-1:17*12]<=12'b111000000000;
			pixels[19*12-1:18*12]<=12'b111000000000;
			pixels[20*12-1:19*12]<=12'b111000000000;
			pixels[21*12-1:20*12]<=12'b111111111111;
			pixels[22*12-1:21*12]<=12'b111111111111;
			pixels[23*12-1:22*12]<=12'b111111111111;
			pixels[24*12-1:23*12]<=12'b111111111111;
		end
		6:begin
			pixels[01*12-1:00*12]<=12'b111111111111;
			pixels[02*12-1:01*12]<=12'b111111111111;
			pixels[03*12-1:02*12]<=12'b111111111111;
			pixels[04*12-1:03*12]<=12'b111111111111;			
			pixels[05*12-1:04*12]<=12'b000000000111;
			pixels[06*12-1:05*12]<=12'b000000000111;
			pixels[07*12-1:06*12]<=12'b000000000111;
			pixels[08*12-1:07*12]<=12'b000000000111;
			pixels[09*12-1:08*12]<=12'b000000000111;
			pixels[10*12-1:09*12]<=12'b000000000111;
			pixels[11*12-1:10*12]<=12'b000000000111;
			pixels[12*12-1:11*12]<=12'b111111111111;
			pixels[13*12-1:12*12]<=12'b111111111111;
			pixels[14*12-1:13*12]<=12'b111000000111;
			pixels[15*12-1:14*12]<=12'b111000000111;
			pixels[16*12-1:15*12]<=12'b111000000111;
			pixels[17*12-1:16*12]<=12'b111000000111;
			pixels[18*12-1:17*12]<=12'b111000000111;
			pixels[19*12-1:18*12]<=12'b111000000111;
			pixels[20*12-1:19*12]<=12'b111000000111;
			pixels[21*12-1:20*12]<=12'b111111111111;
			pixels[22*12-1:21*12]<=12'b111111111111;
			pixels[23*12-1:22*12]<=12'b111111111111;
			pixels[24*12-1:23*12]<=12'b111111111111;
		end
		7:begin
			pixels[01*12-1:00*12]<=12'b111111111111;
			pixels[02*12-1:01*12]<=12'b111111111111;
			pixels[03*12-1:02*12]<=12'b111111111111;
			pixels[04*12-1:03*12]<=12'b111111111111;			
			pixels[05*12-1:04*12]<=12'b111000000111;
			pixels[06*12-1:05*12]<=12'b111000000111;
			pixels[07*12-1:06*12]<=12'b111000000111;
			pixels[08*12-1:07*12]<=12'b111000000111;
			pixels[09*12-1:08*12]<=12'b111000000111;
			pixels[10*12-1:09*12]<=12'b111000000111;
			pixels[11*12-1:10*12]<=12'b111000000111;
			pixels[12*12-1:11*12]<=12'b111000000000;
			pixels[13*12-1:12*12]<=12'b111000000000;
			pixels[14*12-1:13*12]<=12'b111000000000;
			pixels[15*12-1:14*12]<=12'b111000000000;
			pixels[16*12-1:15*12]<=12'b111000000000;
			pixels[17*12-1:16*12]<=12'b111000000000;
			pixels[18*12-1:17*12]<=12'b111000000000;
			pixels[19*12-1:18*12]<=12'b111000000000;
			pixels[20*12-1:19*12]<=12'b111000000000;
			pixels[21*12-1:20*12]<=12'b111000000000;
			pixels[22*12-1:21*12]<=12'b111000000000;
			pixels[23*12-1:22*12]<=12'b111000000000;
			pixels[24*12-1:23*12]<=12'b111000000000;
		end
		8:begin
			pixels[01*12-1:00*12]<=12'b111111111111;
			pixels[02*12-1:01*12]<=12'b111111111111;
			pixels[03*12-1:02*12]<=12'b111111111111;
			pixels[04*12-1:03*12]<=12'b111111111111;			
			pixels[05*12-1:04*12]<=12'b111000000111;
			pixels[06*12-1:05*12]<=12'b111000000111;
			pixels[07*12-1:06*12]<=12'b111000000111;
			pixels[08*12-1:07*12]<=12'b111000000111;
			pixels[09*12-1:08*12]<=12'b111000000111;
			pixels[10*12-1:09*12]<=12'b111000000111;
			pixels[11*12-1:10*12]<=12'b111000000111;
			pixels[12*12-1:11*12]<=12'b111111111111;
			pixels[13*12-1:12*12]<=12'b111111111111;
			pixels[14*12-1:13*12]<=12'b111000000111;
			pixels[15*12-1:14*12]<=12'b111000000111;
			pixels[16*12-1:15*12]<=12'b111000000111;
			pixels[17*12-1:16*12]<=12'b111000000111;
			pixels[18*12-1:17*12]<=12'b111000000111;
			pixels[19*12-1:18*12]<=12'b111000000111;
			pixels[20*12-1:19*12]<=12'b111000000111;
			pixels[21*12-1:20*12]<=12'b111111111111;
			pixels[22*12-1:21*12]<=12'b111111111111;
			pixels[23*12-1:22*12]<=12'b111111111111;
			pixels[24*12-1:23*12]<=12'b111111111111;
		end
		9:begin
			pixels[01*12-1:00*12]<=12'b111111111111;
			pixels[02*12-1:01*12]<=12'b111111111111;
			pixels[03*12-1:02*12]<=12'b111111111111;
			pixels[04*12-1:03*12]<=12'b111111111111;			
			pixels[05*12-1:04*12]<=12'b111000000111;
			pixels[06*12-1:05*12]<=12'b111000000111;
			pixels[07*12-1:06*12]<=12'b111000000111;
			pixels[08*12-1:07*12]<=12'b111000000111;
			pixels[09*12-1:08*12]<=12'b111000000111;
			pixels[10*12-1:09*12]<=12'b111000000111;
			pixels[11*12-1:10*12]<=12'b111000000111;
			pixels[12*12-1:11*12]<=12'b111111111111;
			pixels[13*12-1:12*12]<=12'b111111111111;
			pixels[14*12-1:13*12]<=12'b111000000000;
			pixels[15*12-1:14*12]<=12'b111000000000;
			pixels[16*12-1:15*12]<=12'b111000000000;
			pixels[17*12-1:16*12]<=12'b111000000000;
			pixels[18*12-1:17*12]<=12'b111000000000;
			pixels[19*12-1:18*12]<=12'b111000000000;
			pixels[20*12-1:19*12]<=12'b111000000000;
			pixels[21*12-1:20*12]<=12'b111111111111;
			pixels[22*12-1:21*12]<=12'b111111111111;
			pixels[23*12-1:22*12]<=12'b111111111111;
			pixels[24*12-1:23*12]<=12'b111111111111;
		end

////////////////////////////////////////////////////////////////////////////		
		
		
		10:begin  //A
			pixels[01*12-1:00*12]<=12'b000111111000;
			pixels[02*12-1:01*12]<=12'b001111111100;
			pixels[03*12-1:02*12]<=12'b011111111110;
			pixels[04*12-1:03*12]<=12'b011111111110;			
			pixels[05*12-1:04*12]<=12'b111000000111;
			pixels[06*12-1:05*12]<=12'b111000000111;
			pixels[07*12-1:06*12]<=12'b111000000111;
			pixels[08*12-1:07*12]<=12'b111000000111;
			pixels[09*12-1:08*12]<=12'b111000000111;
			pixels[10*12-1:09*12]<=12'b111000000111;
			pixels[11*12-1:10*12]<=12'b111000000111;
			pixels[12*12-1:11*12]<=12'b111111111111;
			pixels[13*12-1:12*12]<=12'b111111111111;
			pixels[14*12-1:13*12]<=12'b111000000111;
			pixels[15*12-1:14*12]<=12'b111000000111;
			pixels[16*12-1:15*12]<=12'b111000000111;
			pixels[17*12-1:16*12]<=12'b111000000111;
			pixels[18*12-1:17*12]<=12'b111000000111;
			pixels[19*12-1:18*12]<=12'b111000000111;
			pixels[20*12-1:19*12]<=12'b111000000111;
			pixels[21*12-1:20*12]<=12'b111000000111;
			pixels[22*12-1:21*12]<=12'b111000000111;
			pixels[23*12-1:22*12]<=12'b111000000111;
			pixels[24*12-1:23*12]<=12'b111000000111;
		end
		
		11:begin  //B
			pixels[01*12-1:00*12]<=12'b000111111111;
			pixels[02*12-1:01*12]<=12'b001111111111;
			pixels[03*12-1:02*12]<=12'b011111111111;
			pixels[04*12-1:03*12]<=12'b111000000111;			
			pixels[05*12-1:04*12]<=12'b111000000111;
			pixels[06*12-1:05*12]<=12'b111000000111;
			pixels[07*12-1:06*12]<=12'b111000000111;
			pixels[08*12-1:07*12]<=12'b111000000111;
			pixels[09*12-1:08*12]<=12'b111000000111;
			pixels[10*12-1:09*12]<=12'b111000000111;
			pixels[11*12-1:10*12]<=12'b011111111111;
			pixels[12*12-1:11*12]<=12'b001111111111;
			pixels[13*12-1:12*12]<=12'b011111111111;
			pixels[14*12-1:13*12]<=12'b111000000111;
			pixels[15*12-1:14*12]<=12'b111000000111;
			pixels[16*12-1:15*12]<=12'b111000000111;
			pixels[17*12-1:16*12]<=12'b111000000111;
			pixels[18*12-1:17*12]<=12'b111000000111;
			pixels[19*12-1:18*12]<=12'b111000000111;
			pixels[20*12-1:19*12]<=12'b111000000111;
			pixels[21*12-1:20*12]<=12'b111000000111;
			pixels[22*12-1:21*12]<=12'b111111111111;
			pixels[23*12-1:22*12]<=12'b011111111111;
			pixels[24*12-1:23*12]<=12'b001111111111;
		end
		
		12:begin  //C
			pixels[01*12-1:00*12]<=12'b001111111100;
			pixels[02*12-1:01*12]<=12'b011111111110;
			pixels[03*12-1:02*12]<=12'b111111111111;
			pixels[04*12-1:03*12]<=12'b111111111111;			
			pixels[05*12-1:04*12]<=12'b111000000111;
			pixels[06*12-1:05*12]<=12'b111000000111;
			pixels[07*12-1:06*12]<=12'b111000000111;
			pixels[08*12-1:07*12]<=12'b000000000111;
			pixels[09*12-1:08*12]<=12'b000000000111;
			pixels[10*12-1:09*12]<=12'b000000000111;
			pixels[11*12-1:10*12]<=12'b000000000111;
			pixels[12*12-1:11*12]<=12'b000000000111;
			pixels[13*12-1:12*12]<=12'b000000000111;
			pixels[14*12-1:13*12]<=12'b000000000111;
			pixels[15*12-1:14*12]<=12'b000000000111;
			pixels[16*12-1:15*12]<=12'b000000000111;
			pixels[17*12-1:16*12]<=12'b000000000111;
			pixels[18*12-1:17*12]<=12'b000000000111;
			pixels[19*12-1:18*12]<=12'b110000000111;
			pixels[20*12-1:19*12]<=12'b110000000111;
			pixels[21*12-1:20*12]<=12'b111111111111;
			pixels[22*12-1:21*12]<=12'b111111111111;
			pixels[23*12-1:22*12]<=12'b011111111110;
			pixels[24*12-1:23*12]<=12'b001111111100;
		end
		
		13:begin  //D
			pixels[01*12-1:00*12]<=12'b000001111111;
			pixels[02*12-1:01*12]<=12'b000111111111;
			pixels[03*12-1:02*12]<=12'b001111111111;
			pixels[04*12-1:03*12]<=12'b011110000111;
			pixels[05*12-1:04*12]<=12'b011100000111;
			pixels[06*12-1:05*12]<=12'b111000000111;
			pixels[07*12-1:06*12]<=12'b111000000111;
			pixels[08*12-1:07*12]<=12'b111000000111;
			pixels[09*12-1:08*12]<=12'b111000000111;
			pixels[10*12-1:09*12]<=12'b111000000111;
			pixels[11*12-1:10*12]<=12'b111000000111;
			pixels[12*12-1:11*12]<=12'b111000000111;
			pixels[13*12-1:12*12]<=12'b111000000111;
			pixels[14*12-1:13*12]<=12'b111000000111;
			pixels[15*12-1:14*12]<=12'b111000000111;
			pixels[16*12-1:15*12]<=12'b111000000111;
			pixels[17*12-1:16*12]<=12'b111000000111;
			pixels[18*12-1:17*12]<=12'b111000000111;
			pixels[19*12-1:18*12]<=12'b111000000111;
			pixels[20*12-1:19*12]<=12'b111100000111;
			pixels[21*12-1:20*12]<=12'b011110000111;
			pixels[22*12-1:21*12]<=12'b011111111111;
			pixels[23*12-1:22*12]<=12'b001111111111;
			pixels[24*12-1:23*12]<=12'b000011111111;
		end
		
		14:begin  //E
			pixels[01*12-1:00*12]<=12'b111111111111;
			pixels[02*12-1:01*12]<=12'b111111111111;
			pixels[03*12-1:02*12]<=12'b111111111111;
			pixels[04*12-1:03*12]<=12'b110000000111;
			pixels[05*12-1:04*12]<=12'b000000000111;
			pixels[06*12-1:05*12]<=12'b000000000111;
			pixels[07*12-1:06*12]<=12'b000000000111;
			pixels[08*12-1:07*12]<=12'b000000000111;
			pixels[09*12-1:08*12]<=12'b000000000111;
			pixels[10*12-1:09*12]<=12'b000000000111;
			pixels[11*12-1:10*12]<=12'b111111111111;
			pixels[12*12-1:11*12]<=12'b111111111111;
			pixels[13*12-1:12*12]<=12'b111111111111;
			pixels[14*12-1:13*12]<=12'b000000000111;
			pixels[15*12-1:14*12]<=12'b000000000111;
			pixels[16*12-1:15*12]<=12'b000000000111;
			pixels[17*12-1:16*12]<=12'b000000000111;
			pixels[18*12-1:17*12]<=12'b000000000111;
			pixels[19*12-1:18*12]<=12'b000000000111;
			pixels[20*12-1:19*12]<=12'b000000000111;
			pixels[21*12-1:20*12]<=12'b110000000111;
			pixels[22*12-1:21*12]<=12'b111111111111;
			pixels[23*12-1:22*12]<=12'b111111111111;
			pixels[24*12-1:23*12]<=12'b111111111111;
		end
		
		15:begin  //F
			pixels[01*12-1:00*12]<=12'b111111111111;
			pixels[02*12-1:01*12]<=12'b111111111111;
			pixels[03*12-1:02*12]<=12'b111111111111;
			pixels[04*12-1:03*12]<=12'b110000000111;
			pixels[05*12-1:04*12]<=12'b110000000111;
			pixels[06*12-1:05*12]<=12'b000000000111;
			pixels[07*12-1:06*12]<=12'b000000000111;
			pixels[08*12-1:07*12]<=12'b000000000111;
			pixels[09*12-1:08*12]<=12'b000000000111;
			pixels[10*12-1:09*12]<=12'b000000000111;
			pixels[11*12-1:10*12]<=12'b111111111111;
			pixels[12*12-1:11*12]<=12'b111111111111;
			pixels[13*12-1:12*12]<=12'b111111111111;
			pixels[14*12-1:13*12]<=12'b000000000111;
			pixels[15*12-1:14*12]<=12'b000000000111;
			pixels[16*12-1:15*12]<=12'b000000000111;
			pixels[17*12-1:16*12]<=12'b000000000111;
			pixels[18*12-1:17*12]<=12'b000000000111;
			pixels[19*12-1:18*12]<=12'b000000000111;
			pixels[20*12-1:19*12]<=12'b000000000111;
			pixels[21*12-1:20*12]<=12'b000000000111;
			pixels[22*12-1:21*12]<=12'b000000000111;
			pixels[23*12-1:22*12]<=12'b000000000111;
			pixels[24*12-1:23*12]<=12'b000000000111;
		end
		
		16:begin  //G
			pixels[01*12-1:00*12]<=12'b011111111100;
			pixels[02*12-1:01*12]<=12'b111111111110;
			pixels[03*12-1:02*12]<=12'b111111111111;
			pixels[04*12-1:03*12]<=12'b110000001111;
			pixels[05*12-1:04*12]<=12'b000000000111;
			pixels[06*12-1:05*12]<=12'b000000000111;
			pixels[07*12-1:06*12]<=12'b000000000111;
			pixels[08*12-1:07*12]<=12'b000000000111;
			pixels[09*12-1:08*12]<=12'b000000000111;
			pixels[10*12-1:09*12]<=12'b000000000111;
			pixels[11*12-1:10*12]<=12'b000000000111;
			pixels[12*12-1:11*12]<=12'b000000000111;
			pixels[13*12-1:12*12]<=12'b000000000111;
			pixels[14*12-1:13*12]<=12'b111111000111;
			pixels[15*12-1:14*12]<=12'b111111000111;
			pixels[16*12-1:15*12]<=12'b111100000111;
			pixels[17*12-1:16*12]<=12'b110000000111;
			pixels[18*12-1:17*12]<=12'b110000000111;
			pixels[19*12-1:18*12]<=12'b110000000111;
			pixels[20*12-1:19*12]<=12'b110000001111;
			pixels[21*12-1:20*12]<=12'b110000011111;
			pixels[22*12-1:21*12]<=12'b111111111111;
			pixels[23*12-1:22*12]<=12'b011111111110;
			pixels[24*12-1:23*12]<=12'b011111111100;
		end
		
		17:begin  //H
			pixels[01*12-1:00*12]<=12'b111110011111;
			pixels[02*12-1:01*12]<=12'b011100001110;
			pixels[03*12-1:02*12]<=12'b011100001110;
			pixels[04*12-1:03*12]<=12'b011100001110;
			pixels[05*12-1:04*12]<=12'b011100001110;
			pixels[06*12-1:05*12]<=12'b011100001110;
			pixels[07*12-1:06*12]<=12'b011100001110;
			pixels[08*12-1:07*12]<=12'b011100001110;
			pixels[09*12-1:08*12]<=12'b011100001110;
			pixels[10*12-1:09*12]<=12'b011100001110;
			pixels[11*12-1:10*12]<=12'b011111111110;
			pixels[12*12-1:11*12]<=12'b011111111110;
			pixels[13*12-1:12*12]<=12'b011111111110;
			pixels[14*12-1:13*12]<=12'b011111111110;
			pixels[15*12-1:14*12]<=12'b011100001110;
			pixels[16*12-1:15*12]<=12'b011100001110;
			pixels[17*12-1:16*12]<=12'b011100001110;
			pixels[18*12-1:17*12]<=12'b011100001110;
			pixels[19*12-1:18*12]<=12'b011100001110;
			pixels[20*12-1:19*12]<=12'b011100001110;
			pixels[21*12-1:20*12]<=12'b011100001110;
			pixels[22*12-1:21*12]<=12'b011100001110;
			pixels[23*12-1:22*12]<=12'b011100001110;
			pixels[24*12-1:23*12]<=12'b111110011111;
		end
		
		18:begin  //I
			pixels[01*12-1:00*12]<=12'b011111111110;
			pixels[02*12-1:01*12]<=12'b011111111110;
			pixels[03*12-1:02*12]<=12'b000011110000;
			pixels[04*12-1:03*12]<=12'b000011110000;
			pixels[05*12-1:04*12]<=12'b000011110000;
			pixels[06*12-1:05*12]<=12'b000011110000;
			pixels[07*12-1:06*12]<=12'b000011110000;
			pixels[08*12-1:07*12]<=12'b000011110000;
			pixels[09*12-1:08*12]<=12'b000011110000;
			pixels[10*12-1:09*12]<=12'b000011110000;
			pixels[11*12-1:10*12]<=12'b000011110000;
			pixels[12*12-1:11*12]<=12'b000011110000;
			pixels[13*12-1:12*12]<=12'b000011110000;
			pixels[14*12-1:13*12]<=12'b000011110000;
			pixels[15*12-1:14*12]<=12'b000011110000;
			pixels[16*12-1:15*12]<=12'b000011110000;
			pixels[17*12-1:16*12]<=12'b000011110000;
			pixels[18*12-1:17*12]<=12'b000011110000;
			pixels[19*12-1:18*12]<=12'b000011110000;
			pixels[20*12-1:19*12]<=12'b000011110000;
			pixels[21*12-1:20*12]<=12'b000011110000;
			pixels[22*12-1:21*12]<=12'b000011110000;
			pixels[23*12-1:22*12]<=12'b011111111110;
			pixels[24*12-1:23*12]<=12'b011111111110;
		end
		
		19:begin  //J
			pixels[01*12-1:00*12]<=12'b111111111111;
			pixels[02*12-1:01*12]<=12'b111111111111;
			pixels[03*12-1:02*12]<=12'b111111111111;
			pixels[04*12-1:03*12]<=12'b001111000000;
			pixels[05*12-1:04*12]<=12'b001111000000;
			pixels[06*12-1:05*12]<=12'b001111000000;
			pixels[07*12-1:06*12]<=12'b001111000000;
			pixels[08*12-1:07*12]<=12'b001111000000;
			pixels[09*12-1:08*12]<=12'b001111000000;
			pixels[10*12-1:09*12]<=12'b001111000000;
			pixels[11*12-1:10*12]<=12'b001111000000;
			pixels[12*12-1:11*12]<=12'b001111000000;
			pixels[13*12-1:12*12]<=12'b001111000000;
			pixels[14*12-1:13*12]<=12'b001111000000;
			pixels[15*12-1:14*12]<=12'b001111000000;
			pixels[16*12-1:15*12]<=12'b001111000000;
			pixels[17*12-1:16*12]<=12'b001111000000;
			pixels[18*12-1:17*12]<=12'b001111000000;
			pixels[19*12-1:18*12]<=12'b001111000011;
			pixels[20*12-1:19*12]<=12'b001111000011;
			pixels[21*12-1:20*12]<=12'b001111111111;
			pixels[22*12-1:21*12]<=12'b001111111111;
			pixels[23*12-1:22*12]<=12'b000111111110;
			pixels[24*12-1:23*12]<=12'b000011111100;
		end
		
		20:begin  //K
			pixels[01*12-1:00*12]<=12'b111110001111;
			pixels[02*12-1:01*12]<=12'b111100000111;
			pixels[03*12-1:02*12]<=12'b111100000111;
			pixels[04*12-1:03*12]<=12'b011110000111;
			pixels[05*12-1:04*12]<=12'b011111000111;
			pixels[06*12-1:05*12]<=12'b001111100111;
			pixels[07*12-1:06*12]<=12'b000111110111;
			pixels[08*12-1:07*12]<=12'b000011111111;
			pixels[09*12-1:08*12]<=12'b000001111111;
			pixels[10*12-1:09*12]<=12'b000000111111;
			pixels[11*12-1:10*12]<=12'b000000011111;
			pixels[12*12-1:11*12]<=12'b000000001111;
			pixels[13*12-1:12*12]<=12'b000000001111;
			pixels[14*12-1:13*12]<=12'b000000011111;
			pixels[15*12-1:14*12]<=12'b000000111111;
			pixels[16*12-1:15*12]<=12'b000001111111;
			pixels[17*12-1:16*12]<=12'b000011111111;
			pixels[18*12-1:17*12]<=12'b000111110111;
			pixels[19*12-1:18*12]<=12'b001111100111;
			pixels[20*12-1:19*12]<=12'b011111000111;
			pixels[21*12-1:20*12]<=12'b011110000111;
			pixels[22*12-1:21*12]<=12'b111100000111;
			pixels[23*12-1:22*12]<=12'b111100000111;
			pixels[24*12-1:23*12]<=12'b111110001111;
		end
		
		21:begin  //L
			pixels[01*12-1:00*12]<=12'b000000011111;
			pixels[02*12-1:01*12]<=12'b000000001111;
			pixels[03*12-1:02*12]<=12'b000000000111;
			pixels[04*12-1:03*12]<=12'b000000000111;
			pixels[05*12-1:04*12]<=12'b000000000111;
			pixels[06*12-1:05*12]<=12'b000000000111;
			pixels[07*12-1:06*12]<=12'b000000000111;
			pixels[08*12-1:07*12]<=12'b000000000111;
			pixels[09*12-1:08*12]<=12'b000000000111;
			pixels[10*12-1:09*12]<=12'b000000000111;
			pixels[11*12-1:10*12]<=12'b000000000111;
			pixels[12*12-1:11*12]<=12'b000000000111;
			pixels[13*12-1:12*12]<=12'b000000000111;
			pixels[14*12-1:13*12]<=12'b000000000111;
			pixels[15*12-1:14*12]<=12'b000000000111;
			pixels[16*12-1:15*12]<=12'b000000000111;
			pixels[17*12-1:16*12]<=12'b000000000111;
			pixels[18*12-1:17*12]<=12'b000000000111;
			pixels[19*12-1:18*12]<=12'b000000000111;
			pixels[20*12-1:19*12]<=12'b100000000111;
			pixels[21*12-1:20*12]<=12'b110000000111;
			pixels[22*12-1:21*12]<=12'b111111111111;
			pixels[23*12-1:22*12]<=12'b111111111111;
			pixels[24*12-1:23*12]<=12'b111111111111;
		end
		
		22:begin  //M
			pixels[01*12-1:00*12]<=12'b111000000111;
			pixels[02*12-1:01*12]<=12'b111000000111;
			pixels[03*12-1:02*12]<=12'b111100001111;
			pixels[04*12-1:03*12]<=12'b111100001111;
			pixels[05*12-1:04*12]<=12'b111110011111;
			pixels[06*12-1:05*12]<=12'b110110011111;
			pixels[07*12-1:06*12]<=12'b110111111011;
			pixels[08*12-1:07*12]<=12'b110111111011;
			pixels[09*12-1:08*12]<=12'b110111111011;
			pixels[10*12-1:09*12]<=12'b110011110011;
			pixels[11*12-1:10*12]<=12'b110011110011;
			pixels[12*12-1:11*12]<=12'b110001100011;
			pixels[13*12-1:12*12]<=12'b110001100011;
			pixels[14*12-1:13*12]<=12'b110000000011;
			pixels[15*12-1:14*12]<=12'b110000000011;
			pixels[16*12-1:15*12]<=12'b110000000011;
			pixels[17*12-1:16*12]<=12'b110000000011;
			pixels[18*12-1:17*12]<=12'b110000000011;
			pixels[19*12-1:18*12]<=12'b110000000011;
			pixels[20*12-1:19*12]<=12'b110000000011;
			pixels[21*12-1:20*12]<=12'b110000000011;
			pixels[22*12-1:21*12]<=12'b110000000011;
			pixels[23*12-1:22*12]<=12'b110000000011;
			pixels[24*12-1:23*12]<=12'b111000000111;
		end
		
		23:begin  //N
			pixels[01*12-1:00*12]<=12'b110000000111;
			pixels[02*12-1:01*12]<=12'b110000000111;
			pixels[03*12-1:02*12]<=12'b110000001111;
			pixels[04*12-1:03*12]<=12'b110000001111;
			pixels[05*12-1:04*12]<=12'b110000011111;
			pixels[06*12-1:05*12]<=12'b110000011011;
			pixels[07*12-1:06*12]<=12'b110000011011;
			pixels[08*12-1:07*12]<=12'b110000110011;
			pixels[09*12-1:08*12]<=12'b110000110011;
			pixels[10*12-1:09*12]<=12'b110001110011;
			pixels[11*12-1:10*12]<=12'b110001100011;
			pixels[12*12-1:11*12]<=12'b110001100011;
			pixels[13*12-1:12*12]<=12'b110011100011;
			pixels[14*12-1:13*12]<=12'b110011000011;
			pixels[15*12-1:14*12]<=12'b110011000011;
			pixels[16*12-1:15*12]<=12'b110011000011;
			pixels[17*12-1:16*12]<=12'b110110000011;
			pixels[18*12-1:17*12]<=12'b110110000011;
			pixels[19*12-1:18*12]<=12'b110110000011;
			pixels[20*12-1:19*12]<=12'b111100000011;
			pixels[21*12-1:20*12]<=12'b111100000011;
			pixels[22*12-1:21*12]<=12'b111100000011;
			pixels[23*12-1:22*12]<=12'b111000000011;
			pixels[24*12-1:23*12]<=12'b111000000011;
		end
		
		24:begin  //O
			pixels[01*12-1:00*12]<=12'b000111111000;
			pixels[02*12-1:01*12]<=12'b001111111100;
			pixels[03*12-1:02*12]<=12'b011111111110;
			pixels[04*12-1:03*12]<=12'b111111111111;
			pixels[05*12-1:04*12]<=12'b111100001111;
			pixels[06*12-1:05*12]<=12'b111000000111;
			pixels[07*12-1:06*12]<=12'b111000000111;
			pixels[08*12-1:07*12]<=12'b111000000111;
			pixels[09*12-1:08*12]<=12'b111000000111;
			pixels[10*12-1:09*12]<=12'b111000000111;
			pixels[11*12-1:10*12]<=12'b111000000111;
			pixels[12*12-1:11*12]<=12'b111000000111;
			pixels[13*12-1:12*12]<=12'b111000000111;
			pixels[14*12-1:13*12]<=12'b111000000111;
			pixels[15*12-1:14*12]<=12'b111000000111;
			pixels[16*12-1:15*12]<=12'b111000000111;
			pixels[17*12-1:16*12]<=12'b111000000111;
			pixels[18*12-1:17*12]<=12'b111000000111;
			pixels[19*12-1:18*12]<=12'b111000000111;
			pixels[20*12-1:19*12]<=12'b111100001111;
			pixels[21*12-1:20*12]<=12'b111110011111;
			pixels[22*12-1:21*12]<=12'b011111111110;
			pixels[23*12-1:22*12]<=12'b001111111100;
			pixels[24*12-1:23*12]<=12'b000111111000;
		end
		
		
		25:begin  //P
			pixels[01*12-1:00*12]<=12'b000011111111;
			pixels[02*12-1:01*12]<=12'b001111111111;
			pixels[03*12-1:02*12]<=12'b011111111111;
			pixels[04*12-1:03*12]<=12'b111111111111;
			pixels[05*12-1:04*12]<=12'b111100001111;
			pixels[06*12-1:05*12]<=12'b111000000111;
			pixels[07*12-1:06*12]<=12'b111000000111;
			pixels[08*12-1:07*12]<=12'b111000000111;
			pixels[09*12-1:08*12]<=12'b111000000111;
			pixels[10*12-1:09*12]<=12'b111000000111;
			pixels[11*12-1:10*12]<=12'b111100001111;
			pixels[12*12-1:11*12]<=12'b011111111111;
			pixels[13*12-1:12*12]<=12'b001111111111;
			pixels[14*12-1:13*12]<=12'b000111111111;
			pixels[15*12-1:14*12]<=12'b000000000111;
			pixels[16*12-1:15*12]<=12'b000000000111;
			pixels[17*12-1:16*12]<=12'b000000000111;
			pixels[18*12-1:17*12]<=12'b000000000111;
			pixels[19*12-1:18*12]<=12'b000000000111;
			pixels[20*12-1:19*12]<=12'b000000000111;
			pixels[21*12-1:20*12]<=12'b000000000111;
			pixels[22*12-1:21*12]<=12'b000000000111;
			pixels[23*12-1:22*12]<=12'b000000000111;
			pixels[24*12-1:23*12]<=12'b000000000111;
		end
		
		26:begin  //Q
			pixels[01*12-1:00*12]<=12'b000011110000;
			pixels[02*12-1:01*12]<=12'b001111111100;
			pixels[03*12-1:02*12]<=12'b011111111110;
			pixels[04*12-1:03*12]<=12'b011111111110;
			pixels[05*12-1:04*12]<=12'b111100001111;
			pixels[06*12-1:05*12]<=12'b111000000111;
			pixels[07*12-1:06*12]<=12'b111000000111;
			pixels[08*12-1:07*12]<=12'b111000000111;
			pixels[09*12-1:08*12]<=12'b111000000111;
			pixels[10*12-1:09*12]<=12'b111000000111;
			pixels[11*12-1:10*12]<=12'b111000000111;
			pixels[12*12-1:11*12]<=12'b111000000111;
			pixels[13*12-1:12*12]<=12'b111000000111;
			pixels[14*12-1:13*12]<=12'b111000000111;
			pixels[15*12-1:14*12]<=12'b111000000111;
			pixels[16*12-1:15*12]<=12'b111000000111;
			pixels[17*12-1:16*12]<=12'b111000000111;
			pixels[18*12-1:17*12]<=12'b111011000111;
			pixels[19*12-1:18*12]<=12'b111011000111;
			pixels[20*12-1:19*12]<=12'b111110001111;
			pixels[21*12-1:20*12]<=12'b011100011111;
			pixels[22*12-1:21*12]<=12'b011111111110;
			pixels[23*12-1:22*12]<=12'b110111111100;
			pixels[24*12-1:23*12]<=12'b110011111000;
		end
		
		27:begin  //R
			pixels[01*12-1:00*12]<=12'b000011111111;
			pixels[02*12-1:01*12]<=12'b001111111111;
			pixels[03*12-1:02*12]<=12'b011111111111;
			pixels[04*12-1:03*12]<=12'b111111111111;
			pixels[05*12-1:04*12]<=12'b111100001111;
			pixels[06*12-1:05*12]<=12'b111000000111;
			pixels[07*12-1:06*12]<=12'b111000000111;
			pixels[08*12-1:07*12]<=12'b111000000111;
			pixels[09*12-1:08*12]<=12'b111000000111;
			pixels[10*12-1:09*12]<=12'b111000000111;
			pixels[11*12-1:10*12]<=12'b111100001111;
			pixels[12*12-1:11*12]<=12'b011111111111;
			pixels[13*12-1:12*12]<=12'b001111111111;
			pixels[14*12-1:13*12]<=12'b000111111111;
			pixels[15*12-1:14*12]<=12'b000000001111;
			pixels[16*12-1:15*12]<=12'b000000011111;
			pixels[17*12-1:16*12]<=12'b000000111111;
			pixels[18*12-1:17*12]<=12'b000001111111;
			pixels[19*12-1:18*12]<=12'b000011110111;
			pixels[20*12-1:19*12]<=12'b000111100111;
			pixels[21*12-1:20*12]<=12'b001111000111;
			pixels[22*12-1:21*12]<=12'b011110000111;
			pixels[23*12-1:22*12]<=12'b111100000111;
			pixels[24*12-1:23*12]<=12'b111110001111;
		end
		
		28:begin  //S
			pixels[01*12-1:00*12]<=12'b000111111000;
			pixels[02*12-1:01*12]<=12'b011111111110;
			pixels[03*12-1:02*12]<=12'b011111111110;
			pixels[04*12-1:03*12]<=12'b111111111111;
			pixels[05*12-1:04*12]<=12'b111000011111;
			pixels[06*12-1:05*12]<=12'b110000001111;
			pixels[07*12-1:06*12]<=12'b000000000111;
			pixels[08*12-1:07*12]<=12'b000000000111;
			pixels[09*12-1:08*12]<=12'b000000000111;
			pixels[10*12-1:09*12]<=12'b000000001111;
			pixels[11*12-1:10*12]<=12'b000000011111;
			pixels[12*12-1:11*12]<=12'b000111111110;
			pixels[13*12-1:12*12]<=12'b011111111100;
			pixels[14*12-1:13*12]<=12'b011111111000;
			pixels[15*12-1:14*12]<=12'b111110000000;
			pixels[16*12-1:15*12]<=12'b111100000000;
			pixels[17*12-1:16*12]<=12'b111000000000;
			pixels[18*12-1:17*12]<=12'b111000000000;
			pixels[19*12-1:18*12]<=12'b111100000011;
			pixels[20*12-1:19*12]<=12'b111110000111;
			pixels[21*12-1:20*12]<=12'b111111111111;
			pixels[22*12-1:21*12]<=12'b011111111110;
			pixels[23*12-1:22*12]<=12'b011111111110;
			pixels[24*12-1:23*12]<=12'b000111111000;
		end
		
		29:begin  //T
			pixels[01*12-1:00*12]<=12'b111111111111;
			pixels[02*12-1:01*12]<=12'b111111111111;
			pixels[03*12-1:02*12]<=12'b111111111111;
			pixels[04*12-1:03*12]<=12'b000011110000;
			pixels[05*12-1:04*12]<=12'b000011110000;
			pixels[06*12-1:05*12]<=12'b000011110000;
			pixels[07*12-1:06*12]<=12'b000011110000;
			pixels[08*12-1:07*12]<=12'b000011110000;
			pixels[09*12-1:08*12]<=12'b000011110000;
			pixels[10*12-1:09*12]<=12'b000011110000;
			pixels[11*12-1:10*12]<=12'b000011110000;
			pixels[12*12-1:11*12]<=12'b000011110000;
			pixels[13*12-1:12*12]<=12'b000011110000;
			pixels[14*12-1:13*12]<=12'b000011110000;
			pixels[15*12-1:14*12]<=12'b000011110000;
			pixels[16*12-1:15*12]<=12'b000011110000;
			pixels[17*12-1:16*12]<=12'b000011110000;
			pixels[18*12-1:17*12]<=12'b000011110000;
			pixels[19*12-1:18*12]<=12'b000011110000;
			pixels[20*12-1:19*12]<=12'b000011110000;
			pixels[21*12-1:20*12]<=12'b000011110000;
			pixels[22*12-1:21*12]<=12'b000011110000;
			pixels[23*12-1:22*12]<=12'b000011110000;
			pixels[24*12-1:23*12]<=12'b000011110000;
		end
		
		30:begin  //U
			pixels[01*12-1:00*12]<=12'b111110011111;
			pixels[02*12-1:01*12]<=12'b111110011111;
			pixels[03*12-1:02*12]<=12'b011100001110;
			pixels[04*12-1:03*12]<=12'b011100001110;
			pixels[05*12-1:04*12]<=12'b011100001110;
			pixels[06*12-1:05*12]<=12'b011100001110;
			pixels[07*12-1:06*12]<=12'b011100001110;
			pixels[08*12-1:07*12]<=12'b011100001110;
			pixels[09*12-1:08*12]<=12'b011100001110;
			pixels[10*12-1:09*12]<=12'b011100001110;
			pixels[11*12-1:10*12]<=12'b011100001110;
			pixels[12*12-1:11*12]<=12'b011100001110;
			pixels[13*12-1:12*12]<=12'b011100001110;
			pixels[14*12-1:13*12]<=12'b011100001110;
			pixels[15*12-1:14*12]<=12'b011100001110;
			pixels[16*12-1:15*12]<=12'b011100001110;
			pixels[17*12-1:16*12]<=12'b011100001110;
			pixels[18*12-1:17*12]<=12'b011100001110;
			pixels[19*12-1:18*12]<=12'b011100001110;
			pixels[20*12-1:19*12]<=12'b011100001110;
			pixels[21*12-1:20*12]<=12'b011110011110;
			pixels[22*12-1:21*12]<=12'b011111111110;
			pixels[23*12-1:22*12]<=12'b001111111100;
			pixels[24*12-1:23*12]<=12'b000111111000;
		end
		
		31:begin  //V
			pixels[01*12-1:00*12]<=12'b111000000111;
			pixels[02*12-1:01*12]<=12'b111000000111;
			pixels[03*12-1:02*12]<=12'b111000000111;
			pixels[04*12-1:03*12]<=12'b111000000111;
			pixels[05*12-1:04*12]<=12'b111000000111;
			pixels[06*12-1:05*12]<=12'b111000000111;
			pixels[07*12-1:06*12]<=12'b111000000111;
			pixels[08*12-1:07*12]<=12'b111000000111;
			pixels[09*12-1:08*12]<=12'b111000000111;
			pixels[10*12-1:09*12]<=12'b011100001110;
			pixels[11*12-1:10*12]<=12'b011100001110;
			pixels[12*12-1:11*12]<=12'b011100001110;
			pixels[13*12-1:12*12]<=12'b011100001110;
			pixels[14*12-1:13*12]<=12'b011100001110;
			pixels[15*12-1:14*12]<=12'b011100001110;
			pixels[16*12-1:15*12]<=12'b011100001110;
			pixels[17*12-1:16*12]<=12'b001110011100;
			pixels[18*12-1:17*12]<=12'b001110011100;
			pixels[19*12-1:18*12]<=12'b001110011100;
			pixels[20*12-1:19*12]<=12'b001111111100;
			pixels[21*12-1:20*12]<=12'b000111111000;
			pixels[22*12-1:21*12]<=12'b000111111000;
			pixels[23*12-1:22*12]<=12'b000011110000;
			pixels[24*12-1:23*12]<=12'b000011110000;
		end
		
		32:begin  //W
			pixels[01*12-1:00*12]<=12'b111000000111;
			pixels[02*12-1:01*12]<=12'b110000000011;
			pixels[03*12-1:02*12]<=12'b110000000011;
			pixels[04*12-1:03*12]<=12'b110000000011;
			pixels[05*12-1:04*12]<=12'b110000000011;
			pixels[06*12-1:05*12]<=12'b110000000011;
			pixels[07*12-1:06*12]<=12'b110000000011;
			pixels[08*12-1:07*12]<=12'b110000000011;
			pixels[09*12-1:08*12]<=12'b110000000011;
			pixels[10*12-1:09*12]<=12'b110001100011;
			pixels[11*12-1:10*12]<=12'b110001100011;
			pixels[12*12-1:11*12]<=12'b110001100011;
			pixels[13*12-1:12*12]<=12'b110011110011;
			pixels[14*12-1:13*12]<=12'b110011110011;
			pixels[15*12-1:14*12]<=12'b110011111011;
			pixels[16*12-1:15*12]<=12'b110111111011;
			pixels[17*12-1:16*12]<=12'b111111111111;
			pixels[18*12-1:17*12]<=12'b111111111111;
			pixels[19*12-1:18*12]<=12'b111110011111;
			pixels[20*12-1:19*12]<=12'b111110011111;
			pixels[21*12-1:20*12]<=12'b111100001111;
			pixels[22*12-1:21*12]<=12'b111100001111;
			pixels[23*12-1:22*12]<=12'b111000000111;
			pixels[24*12-1:23*12]<=12'b111000000111;
		end
		
		33:begin  //X
			pixels[01*12-1:00*12]<=12'b111000000111;
			pixels[02*12-1:01*12]<=12'b111000000111;
			pixels[03*12-1:02*12]<=12'b111100001111;
			pixels[04*12-1:03*12]<=12'b011100001110;
			pixels[05*12-1:04*12]<=12'b011100001110;
			pixels[06*12-1:05*12]<=12'b001110011100;
			pixels[07*12-1:06*12]<=12'b001110011100;
			pixels[08*12-1:07*12]<=12'b001110011100;
			pixels[09*12-1:08*12]<=12'b000110011000;
			pixels[10*12-1:09*12]<=12'b000111111000;
			pixels[11*12-1:10*12]<=12'b000011110000;
			pixels[12*12-1:11*12]<=12'b000011110000;
			pixels[13*12-1:12*12]<=12'b000011110000;
			pixels[14*12-1:13*12]<=12'b000011110000;
			pixels[15*12-1:14*12]<=12'b000111111000;
			pixels[16*12-1:15*12]<=12'b000111111000;
			pixels[17*12-1:16*12]<=12'b001111111100;
			pixels[18*12-1:17*12]<=12'b001110011100;
			pixels[19*12-1:18*12]<=12'b001110011100;
			pixels[20*12-1:19*12]<=12'b011110011110;
			pixels[21*12-1:20*12]<=12'b011100001110;
			pixels[22*12-1:21*12]<=12'b111000000111;
			pixels[23*12-1:22*12]<=12'b111000000111;
			pixels[24*12-1:23*12]<=12'b111000000111;
		end
		
		34:begin  //Y
			pixels[01*12-1:00*12]<=12'b111000000111;
			pixels[02*12-1:01*12]<=12'b111000000111;
			pixels[03*12-1:02*12]<=12'b111000000111;
			pixels[04*12-1:03*12]<=12'b111000000111;
			pixels[05*12-1:04*12]<=12'b111100001111;
			pixels[06*12-1:05*12]<=12'b011100001110;
			pixels[07*12-1:06*12]<=12'b011100001110;
			pixels[08*12-1:07*12]<=12'b001110011100;
			pixels[09*12-1:08*12]<=12'b001110011100;
			pixels[10*12-1:09*12]<=12'b001111111100;
			pixels[11*12-1:10*12]<=12'b000111111000;
			pixels[12*12-1:11*12]<=12'b000111111000;
			pixels[13*12-1:12*12]<=12'b000111111000;
			pixels[14*12-1:13*12]<=12'b000011110000;
			pixels[15*12-1:14*12]<=12'b000011110000;
			pixels[16*12-1:15*12]<=12'b000011110000;
			pixels[17*12-1:16*12]<=12'b000011110000;
			pixels[18*12-1:17*12]<=12'b000011110000;
			pixels[19*12-1:18*12]<=12'b000011110000;
			pixels[20*12-1:19*12]<=12'b000011110000;
			pixels[21*12-1:20*12]<=12'b000011110000;
			pixels[22*12-1:21*12]<=12'b000011110000;
			pixels[23*12-1:22*12]<=12'b000011110000;
			pixels[24*12-1:23*12]<=12'b000011110000;
		end
		
		35:begin  //Z
			pixels[01*12-1:00*12]<=12'b111111111111;
			pixels[02*12-1:01*12]<=12'b111111111111;
			pixels[03*12-1:02*12]<=12'b111111111111;
			pixels[04*12-1:03*12]<=12'b111000000000;
			pixels[05*12-1:04*12]<=12'b011100000000;
			pixels[06*12-1:05*12]<=12'b011100000000;
			pixels[07*12-1:06*12]<=12'b001110000000;
			pixels[08*12-1:07*12]<=12'b001110000000;
			pixels[09*12-1:08*12]<=12'b000111000000;
			pixels[10*12-1:09*12]<=12'b000111000000;
			pixels[11*12-1:10*12]<=12'b000011100000;
			pixels[12*12-1:11*12]<=12'b000011100000;
			pixels[13*12-1:12*12]<=12'b000001110000;
			pixels[14*12-1:13*12]<=12'b000001110000;
			pixels[15*12-1:14*12]<=12'b000000111000;
			pixels[16*12-1:15*12]<=12'b000000111000;
			pixels[17*12-1:16*12]<=12'b000000011100;
			pixels[18*12-1:17*12]<=12'b000000011100;
			pixels[19*12-1:18*12]<=12'b000000001110;
			pixels[20*12-1:19*12]<=12'b000000001110;
			pixels[21*12-1:20*12]<=12'b000000000111;
			pixels[22*12-1:21*12]<=12'b111111111111;
			pixels[23*12-1:22*12]<=12'b111111111111;
			pixels[24*12-1:23*12]<=12'b111111111111;
		end
		
		36:begin  //:
			pixels[01*12-1:00*12]<=12'b000000000000;
			pixels[02*12-1:01*12]<=12'b000000000000;
			pixels[03*12-1:02*12]<=12'b000000000000;
			pixels[04*12-1:03*12]<=12'b000000000000;
			pixels[05*12-1:04*12]<=12'b000001100000;
			pixels[06*12-1:05*12]<=12'b000011110000;
			pixels[07*12-1:06*12]<=12'b000011110000;
			pixels[08*12-1:07*12]<=12'b000011110000;
			pixels[09*12-1:08*12]<=12'b000001100000;
			pixels[10*12-1:09*12]<=12'b000000000000;
			pixels[11*12-1:10*12]<=12'b000000000000;
			pixels[12*12-1:11*12]<=12'b000000000000;
			pixels[13*12-1:12*12]<=12'b000000000000;
			pixels[14*12-1:13*12]<=12'b000000000000;
			pixels[15*12-1:14*12]<=12'b000000000000;
			pixels[16*12-1:15*12]<=12'b000001100000;
			pixels[17*12-1:16*12]<=12'b000011110000;
			pixels[18*12-1:17*12]<=12'b000011110000;
			pixels[19*12-1:18*12]<=12'b000011110000;
			pixels[20*12-1:19*12]<=12'b000001100000;
			pixels[21*12-1:20*12]<=12'b000000000000;
			pixels[22*12-1:21*12]<=12'b000000000000;
			pixels[23*12-1:22*12]<=12'b000000000000;
			pixels[24*12-1:23*12]<=12'b000000000000;
		end
		
		37:begin  //▲
			pixels[01*12-1:00*12]<=12'b000000000000;
			pixels[02*12-1:01*12]<=12'b000000000000;
			pixels[03*12-1:02*12]<=12'b000000000000;
			pixels[04*12-1:03*12]<=12'b000000000000;
			pixels[05*12-1:04*12]<=12'b000000000000;
			pixels[06*12-1:05*12]<=12'b000000000000;
			pixels[07*12-1:06*12]<=12'b000000000000;
			pixels[08*12-1:07*12]<=12'b000000000000;
			pixels[09*12-1:08*12]<=12'b000000000000;
			pixels[10*12-1:09*12]<=12'b000001100000;
			pixels[11*12-1:10*12]<=12'b000011110000;
			pixels[12*12-1:11*12]<=12'b000111111000;
			pixels[13*12-1:12*12]<=12'b001111111100;
			pixels[14*12-1:13*12]<=12'b011111111110;
			pixels[15*12-1:14*12]<=12'b111111111111;
			pixels[16*12-1:15*12]<=12'b111111111111;
			pixels[17*12-1:16*12]<=12'b000000000000;
			pixels[18*12-1:17*12]<=12'b000000000000;
			pixels[19*12-1:18*12]<=12'b000000000000;
			pixels[20*12-1:19*12]<=12'b000000000000;
			pixels[21*12-1:20*12]<=12'b000000000000;
			pixels[22*12-1:21*12]<=12'b000000000000;
			pixels[23*12-1:22*12]<=12'b000000000000;
			pixels[24*12-1:23*12]<=12'b000000000000;
		end
		
		38:begin  //▼
			pixels[01*12-1:00*12]<=12'b000000000000;
			pixels[02*12-1:01*12]<=12'b000000000000;
			pixels[03*12-1:02*12]<=12'b000000000000;
			pixels[04*12-1:03*12]<=12'b000000000000;
			pixels[05*12-1:04*12]<=12'b000000000000;
			pixels[06*12-1:05*12]<=12'b000000000000;
			pixels[07*12-1:06*12]<=12'b000000000000;
			pixels[08*12-1:07*12]<=12'b000000000000;
			pixels[09*12-1:08*12]<=12'b000000000000;
			pixels[10*12-1:09*12]<=12'b111111111111;
			pixels[11*12-1:10*12]<=12'b111111111111;
			pixels[12*12-1:11*12]<=12'b011111111110;
			pixels[13*12-1:12*12]<=12'b001111111100;
			pixels[14*12-1:13*12]<=12'b000111111000;
			pixels[15*12-1:14*12]<=12'b000011110000;
			pixels[16*12-1:15*12]<=12'b000001100000;
			pixels[17*12-1:16*12]<=12'b000000000000;
			pixels[18*12-1:17*12]<=12'b000000000000;
			pixels[19*12-1:18*12]<=12'b000000000000;
			pixels[20*12-1:19*12]<=12'b000000000000;
			pixels[21*12-1:20*12]<=12'b000000000000;
			pixels[22*12-1:21*12]<=12'b000000000000;
			pixels[23*12-1:22*12]<=12'b000000000000;
			pixels[24*12-1:23*12]<=12'b000000000000;
			
		end
		
		39:begin  //^
			pixels[01*12-1:00*12]<=12'b000000000000;
			pixels[02*12-1:01*12]<=12'b000000000000;
			pixels[03*12-1:02*12]<=12'b000000000000;
			pixels[04*12-1:03*12]<=12'b000000000000;
			pixels[05*12-1:04*12]<=12'b000000000000;
			pixels[06*12-1:05*12]<=12'b000000000000;
			pixels[07*12-1:06*12]<=12'b000000000000;
			pixels[08*12-1:07*12]<=12'b000000000000;
			pixels[09*12-1:08*12]<=12'b000000000000;
			pixels[10*12-1:09*12]<=12'b000001100000;
			pixels[11*12-1:10*12]<=12'b000011110000;
			pixels[12*12-1:11*12]<=12'b000110011000;
			pixels[13*12-1:12*12]<=12'b001100001100;
			pixels[14*12-1:13*12]<=12'b011000000110;
			pixels[15*12-1:14*12]<=12'b110000000011;
			pixels[16*12-1:15*12]<=12'b100000000001;
			pixels[17*12-1:16*12]<=12'b000000000000;
			pixels[18*12-1:17*12]<=12'b000000000000;
			pixels[19*12-1:18*12]<=12'b000000000000;
			pixels[20*12-1:19*12]<=12'b000000000000;
			pixels[21*12-1:20*12]<=12'b000000000000;
			pixels[22*12-1:21*12]<=12'b000000000000;
			pixels[23*12-1:22*12]<=12'b000000000000;
			pixels[24*12-1:23*12]<=12'b000000000000;
		end
		
		40:begin  //ˇ
			pixels[01*12-1:00*12]<=12'b000000000000;
			pixels[02*12-1:01*12]<=12'b000000000000;
			pixels[03*12-1:02*12]<=12'b000000000000;
			pixels[04*12-1:03*12]<=12'b000000000000;
			pixels[05*12-1:04*12]<=12'b000000000000;
			pixels[06*12-1:05*12]<=12'b000000000000;
			pixels[07*12-1:06*12]<=12'b000000000000;
			pixels[08*12-1:07*12]<=12'b000000000000;
			pixels[09*12-1:08*12]<=12'b100000000001;
			pixels[10*12-1:09*12]<=12'b110000000011;
			pixels[11*12-1:10*12]<=12'b011000000110;
			pixels[12*12-1:11*12]<=12'b001100001100;
			pixels[13*12-1:12*12]<=12'b000110011000;
			pixels[14*12-1:13*12]<=12'b000011110000;
			pixels[15*12-1:14*12]<=12'b000001100000;
			pixels[16*12-1:15*12]<=12'b000000000000;
			pixels[17*12-1:16*12]<=12'b000000000000;
			pixels[18*12-1:17*12]<=12'b000000000000;
			pixels[19*12-1:18*12]<=12'b000000000000;
			pixels[20*12-1:19*12]<=12'b000000000000;
			pixels[21*12-1:20*12]<=12'b000000000000;
			pixels[22*12-1:21*12]<=12'b000000000000;
			pixels[23*12-1:22*12]<=12'b000000000000;
			pixels[24*12-1:23*12]<=12'b000000000000;
		end

		
		default:begin
			pixels[12*24-1:0]<=288'b0;
		end
		endcase
		
	end
endmodule